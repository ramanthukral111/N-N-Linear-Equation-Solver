-- LU_Linear_Equation_Solver_tb.vhd

-- Generated using ACDS version 18.1 625

library IEEE;
use IEEE.std_logic_1164.all;
use IEEE.numeric_std.all;

entity LU_Linear_Equation_Solver_tb is
end entity LU_Linear_Equation_Solver_tb;

architecture rtl of LU_Linear_Equation_Solver_tb is
	component LU_Linear_Equation_Solver is
		port (
			clk_clk       : in std_logic := 'X'; -- clk
			reset_reset_n : in std_logic := 'X'  -- reset_n
		);
	end component LU_Linear_Equation_Solver;

	component altera_avalon_clock_source is
		generic (
			CLOCK_RATE : positive := 10;
			CLOCK_UNIT : positive := 1000000
		);
		port (
			clk : out std_logic   -- clk
		);
	end component altera_avalon_clock_source;

	component altera_avalon_reset_source is
		generic (
			ASSERT_HIGH_RESET    : integer := 1;
			INITIAL_RESET_CYCLES : integer := 0
		);
		port (
			reset : out std_logic;        -- reset_n
			clk   : in  std_logic := 'X'  -- clk
		);
	end component altera_avalon_reset_source;

	signal lu_linear_equation_solver_inst_clk_bfm_clk_clk       : std_logic; -- LU_Linear_Equation_Solver_inst_clk_bfm:clk -> [LU_Linear_Equation_Solver_inst:clk_clk, LU_Linear_Equation_Solver_inst_reset_bfm:clk]
	signal lu_linear_equation_solver_inst_reset_bfm_reset_reset : std_logic; -- LU_Linear_Equation_Solver_inst_reset_bfm:reset -> LU_Linear_Equation_Solver_inst:reset_reset_n

begin

	lu_linear_equation_solver_inst : component LU_Linear_Equation_Solver
		port map (
			clk_clk       => lu_linear_equation_solver_inst_clk_bfm_clk_clk,       --   clk.clk
			reset_reset_n => lu_linear_equation_solver_inst_reset_bfm_reset_reset  -- reset.reset_n
		);

	lu_linear_equation_solver_inst_clk_bfm : component altera_avalon_clock_source
		generic map (
			CLOCK_RATE => 50000000,
			CLOCK_UNIT => 1
		)
		port map (
			clk => lu_linear_equation_solver_inst_clk_bfm_clk_clk  -- clk.clk
		);

	lu_linear_equation_solver_inst_reset_bfm : component altera_avalon_reset_source
		generic map (
			ASSERT_HIGH_RESET    => 0,
			INITIAL_RESET_CYCLES => 50
		)
		port map (
			reset => lu_linear_equation_solver_inst_reset_bfm_reset_reset, -- reset.reset_n
			clk   => lu_linear_equation_solver_inst_clk_bfm_clk_clk        --   clk.clk
		);

end architecture rtl; -- of LU_Linear_Equation_Solver_tb
