Float_32_Add_inst : Float_32_Add PORT MAP (
		add_sub	 => add_sub_sig,
		clock	 => clock_sig,
		dataa	 => dataa_sig,
		datab	 => datab_sig,
		result	 => result_sig
	);
