-- megafunction wizard: %ALTFP_DIV%
-- GENERATION: STANDARD
-- VERSION: WM1.0
-- MODULE: altfp_div 

-- ============================================================
-- File Name: Float_32_Div.vhd
-- Megafunction Name(s):
-- 			altfp_div
--
-- Simulation Library Files(s):
-- 			lpm
-- ============================================================
-- ************************************************************
-- THIS IS A WIZARD-GENERATED FILE. DO NOT EDIT THIS FILE!
--
-- 18.1.0 Build 625 09/12/2018 SJ Lite Edition
-- ************************************************************


--Copyright (C) 2018  Intel Corporation. All rights reserved.
--Your use of Intel Corporation's design tools, logic functions 
--and other software and tools, and its AMPP partner logic 
--functions, and any output files from any of the foregoing 
--(including device programming or simulation files), and any 
--associated documentation or information are expressly subject 
--to the terms and conditions of the Intel Program License 
--Subscription Agreement, the Intel Quartus Prime License Agreement,
--the Intel FPGA IP License Agreement, or other applicable license
--agreement, including, without limitation, that your use is for
--the sole purpose of programming logic devices manufactured by
--Intel and sold by Intel or its authorized distributors.  Please
--refer to the applicable agreement for further details.


--altfp_div CBX_AUTO_BLACKBOX="ALL" DENORMAL_SUPPORT="NO" DEVICE_FAMILY="Cyclone IV E" OPTIMIZE="AREA" PIPELINE=33 REDUCED_FUNCTIONALITY="NO" WIDTH_EXP=8 WIDTH_MAN=23 clock dataa datab division_by_zero result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END


--altfp_div_csa CARRY_SELECT="YES" CBX_AUTO_BLACKBOX="ALL" DATAB_IS_CONSTANT="YES" LPM_DIRECTION="ADD" LPM_WIDTH=24 cin cout dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 2 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_csa_gvc IS 
	 PORT 
	 ( 
		 cin	:	IN  STD_LOGIC := '0';
		 cout	:	OUT  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_csa_gvc;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_csa_gvc IS

	 SIGNAL  wire_csa_lower_w_lg_w_lg_cout819w820w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout818w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_cout819w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_csa_lower_w_lg_w_lg_w_lg_cout819w820w821w	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_csa_lower_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_lower_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  wire_vcc	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_cout	:	STD_LOGIC;
	 SIGNAL  wire_csa_upper1_result	:	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  adder_upper_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  cout_w :	STD_LOGIC;
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	wire_vcc <= '1';
	adder_upper_w <= dataa(23 DOWNTO 12);
	cout <= cout_w;
	cout_w <= (wire_csa_lower_cout AND wire_csa_upper1_cout);
	result <= result_w;
	result_w <= ( wire_csa_lower_w_lg_w_lg_w_lg_cout819w820w821w & wire_csa_lower_result);
	loop0 : FOR i IN 0 TO 11 GENERATE 
		wire_csa_lower_w_lg_w_lg_cout819w820w(i) <= wire_csa_lower_w_lg_cout819w(0) AND adder_upper_w(i);
	END GENERATE loop0;
	loop1 : FOR i IN 0 TO 11 GENERATE 
		wire_csa_lower_w_lg_cout818w(i) <= wire_csa_lower_cout AND wire_csa_upper1_result(i);
	END GENERATE loop1;
	wire_csa_lower_w_lg_cout819w(0) <= NOT wire_csa_lower_cout;
	loop2 : FOR i IN 0 TO 11 GENERATE 
		wire_csa_lower_w_lg_w_lg_w_lg_cout819w820w821w(i) <= wire_csa_lower_w_lg_w_lg_cout819w820w(i) OR wire_csa_lower_w_lg_cout818w(i);
	END GENERATE loop2;
	csa_lower :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		cin => cin,
		cout => wire_csa_lower_cout,
		dataa => dataa(11 DOWNTO 0),
		datab => datab(11 DOWNTO 0),
		result => wire_csa_lower_result
	  );
	csa_upper1 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 12
	  )
	  PORT MAP ( 
		cin => wire_vcc,
		cout => wire_csa_upper1_cout,
		dataa => dataa(23 DOWNTO 12),
		datab => datab(23 DOWNTO 12),
		result => wire_csa_upper1_result
	  );

 END RTL; --Float_32_Div_altfp_div_csa_gvc


--altfp_div_srt_ext CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" ITERATION=14 OPTMIZE="AREA" WIDTH_DIV=24 aclr clken clock denom divider numer quotient remain
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END


--altfp_div_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DATAB_IS_CONSTANT="NO" LPM_DIRECTION="ADD" LPM_WIDTH=24 dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_csa_jub IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_csa_jub;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_csa_jub IS

	 SIGNAL  wire_add_sub28_result	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub28_result;
	add_sub28 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 24
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub28_result
	  );

 END RTL; --Float_32_Div_altfp_div_csa_jub


--altfp_div_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DATAB_IS_CONSTANT="NO" LPM_DIRECTION="SUB" LPM_PIPELINE=1 LPM_WIDTH=28 aclr clken clock dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_csa_vse IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 dataa	:	IN  STD_LOGIC_VECTOR (27 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (27 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (27 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_csa_vse;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_csa_vse IS

	 SIGNAL  wire_add_sub29_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub29_result;
	add_sub29 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 28
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub29_result
	  );

 END RTL; --Float_32_Div_altfp_div_csa_vse


--altfp_div_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DATAB_IS_CONSTANT="NO" LPM_DIRECTION="SUB" LPM_WIDTH=28 dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_csa_ovb IS 
	 PORT 
	 ( 
		 dataa	:	IN  STD_LOGIC_VECTOR (27 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (27 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (27 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_csa_ovb;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_csa_ovb IS

	 SIGNAL  wire_add_sub30_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub30_result;
	add_sub30 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 28
	  )
	  PORT MAP ( 
		dataa => dataa,
		datab => datab,
		result => wire_add_sub30_result
	  );

 END RTL; --Float_32_Div_altfp_div_csa_ovb


--srt_block_int CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" OPTIMIZE="AREA" POSITION="FIRST" WIDTH_DIV=24 WIDTH_RK_IN=24 WIDTH_RK_OUT=25 WIDTH_ROM=3 WIDTH_ROM_ADD=12 aclr clken clock divider divider_reg Rk Rk_next rom
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END


--altfp_div_csa CARRY_SELECT="NO" CBX_AUTO_BLACKBOX="ALL" DATAB_IS_CONSTANT="NO" LPM_WIDTH=27 add_sub dataa datab result
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 1 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_csa_lsa IS 
	 PORT 
	 ( 
		 add_sub	:	IN  STD_LOGIC := '1';
		 dataa	:	IN  STD_LOGIC_VECTOR (26 DOWNTO 0) := (OTHERS => '0');
		 datab	:	IN  STD_LOGIC_VECTOR (26 DOWNTO 0) := (OTHERS => '0');
		 result	:	OUT  STD_LOGIC_VECTOR (26 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_csa_lsa;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_csa_lsa IS

	 SIGNAL  wire_add_sub34_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  result_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	result <= result_w;
	result_w <= wire_add_sub34_result;
	add_sub34 :  lpm_add_sub
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 27
	  )
	  PORT MAP ( 
		add_sub => add_sub,
		dataa => dataa,
		datab => datab,
		result => wire_add_sub34_result
	  );

 END RTL; --Float_32_Div_altfp_div_csa_lsa


--qds_block CBX_AUTO_BLACKBOX="ALL" FIRST_QDS="YES" aclr clken clock decoder_bus decoder_output
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_compare 4 lpm_mux 1 reg 2 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_qds_block_7o8 IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 decoder_bus	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
		 decoder_output	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END Float_32_Div_qds_block_7o8;

 ARCHITECTURE RTL OF Float_32_Div_qds_block_7o8 IS

	 SIGNAL	 q_next_dffe	:	STD_LOGIC_VECTOR(1 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr36_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr37_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr38_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr39_aleb	:	STD_LOGIC;
	 SIGNAL  wire_mux35_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_mux35_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_k_comp_w_range1602w1611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_k_comp_w_range1604w1613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_k_comp_w_range1600w1610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_k_comp_w_range1603w1612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_k_comp_w_range1604w1607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1613w1614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1607w1608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  decoder_output_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  Div_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  k_comp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  mk_bus_const_w :	STD_LOGIC_VECTOR (511 DOWNTO 0);
	 SIGNAL  mk_bus_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mk_neg1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos0_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos2_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  q_next_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  Rk_in_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Rk_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_k_comp_w_range1600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_k_comp_w_range1602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_k_comp_w_range1603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_k_comp_w_range1604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block31_w_q_next_w_range1617w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_qds_block31_w_lg_w_k_comp_w_range1602w1611w(0) <= wire_qds_block31_w_k_comp_w_range1602w(0) AND wire_qds_block31_w_lg_w_k_comp_w_range1600w1610w(0);
	wire_qds_block31_w_lg_w_k_comp_w_range1604w1613w(0) <= wire_qds_block31_w_k_comp_w_range1604w(0) AND wire_qds_block31_w_lg_w_k_comp_w_range1603w1612w(0);
	wire_qds_block31_w_lg_w_k_comp_w_range1600w1610w(0) <= NOT wire_qds_block31_w_k_comp_w_range1600w(0);
	wire_qds_block31_w_lg_w_k_comp_w_range1603w1612w(0) <= NOT wire_qds_block31_w_k_comp_w_range1603w(0);
	wire_qds_block31_w_lg_w_k_comp_w_range1604w1607w(0) <= NOT wire_qds_block31_w_k_comp_w_range1604w(0);
	wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1613w1614w(0) <= wire_qds_block31_w_lg_w_k_comp_w_range1604w1613w(0) OR wire_qds_block31_w_lg_w_k_comp_w_range1602w1611w(0);
	wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1607w1608w(0) <= wire_qds_block31_w_lg_w_k_comp_w_range1604w1607w(0) OR wire_qds_block31_w_k_comp_w_range1600w(0);
	decoder_output <= decoder_output_w;
	decoder_output_w <= ( "0" & q_next_dffe);
	Div_w <= decoder_bus(3 DOWNTO 0);
	k_comp_w <= ( wire_cmpr39_aleb & wire_cmpr38_aleb & wire_cmpr37_aleb & wire_cmpr36_aleb);
	mk_bus_const_w <= ( "01011101000111111110000110100011" & "01011010000111101110001010100110" & "01010111000111011110001110101001" & "01010100000111001110010010101100" & "01010001000110111110010110101111" & "01001110000110101110011010110010" & "01001011000110011110011110110101" & "01001000000110001110100010111000" & "01000101000101111110100110111011" & "01000010000101101110101010111110" & "00111111000101011110101111000001" & "00111100000101001110110011000100" & "00111001000100111110110111000111" & "00110110000100101110111011001010" & "00110011000100011110111111001101" & "00110000000100001111000011010000");
	mk_bus_w <= wire_mux35_result;
	mk_neg1_w <= ( mk_bus_w(7) & mk_bus_w(7 DOWNTO 0));
	mk_pos0_w <= ( mk_bus_w(15) & mk_bus_w(15 DOWNTO 8));
	mk_pos1_w <= ( mk_bus_w(23) & mk_bus_w(23 DOWNTO 16));
	mk_pos2_w <= ( mk_bus_w(31) & mk_bus_w(31 DOWNTO 24));
	q_next_w <= ( k_comp_w(1) & wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1607w1608w & wire_qds_block31_w_lg_w_lg_w_k_comp_w_range1604w1613w1614w);
	Rk_in_w <= ( decoder_bus(11 DOWNTO 4) & "0");
	Rk_w <= Rk_in_w;
	wire_qds_block31_w_k_comp_w_range1600w(0) <= k_comp_w(0);
	wire_qds_block31_w_k_comp_w_range1602w(0) <= k_comp_w(1);
	wire_qds_block31_w_k_comp_w_range1603w(0) <= k_comp_w(2);
	wire_qds_block31_w_k_comp_w_range1604w(0) <= k_comp_w(3);
	wire_qds_block31_w_q_next_w_range1617w <= q_next_w(1 DOWNTO 0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_next_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_next_dffe <= wire_qds_block31_w_q_next_w_range1617w;
			END IF;
		END IF;
	END PROCESS;
	cmpr36 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr36_aleb,
		dataa => Rk_w,
		datab => mk_neg1_w
	  );
	cmpr37 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr37_aleb,
		dataa => Rk_w,
		datab => mk_pos0_w
	  );
	cmpr38 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr38_aleb,
		dataa => Rk_w,
		datab => mk_pos1_w
	  );
	cmpr39 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr39_aleb,
		dataa => Rk_w,
		datab => mk_pos2_w
	  );
	loop3 : FOR i IN 0 TO 15 GENERATE
		loop4 : FOR j IN 0 TO 31 GENERATE
			wire_mux35_data_2d(i, j) <= mk_bus_const_w(i*32+j);
		END GENERATE loop4;
	END GENERATE loop3;
	mux35 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_mux35_data_2d,
		result => wire_mux35_result,
		sel => Div_w
	  );

 END RTL; --Float_32_Div_qds_block_7o8

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 1 lpm_compare 4 lpm_mux 2 reg 100 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_srt_block_int_sfk IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 divider	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 divider_reg	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 Rk	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 Rk_next	:	OUT  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 rom	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END Float_32_Div_srt_block_int_sfk;

 ARCHITECTURE RTL OF Float_32_Div_srt_block_int_sfk IS

	 SIGNAL  wire_altfp_div_csa33_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL	 divider_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divider_dffe_1a	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_dffe	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_next_dffe	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_out_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mux32_data_2d	:	STD_LOGIC_2D(3 DOWNTO 0, 26 DOWNTO 0);
	 SIGNAL  wire_mux32_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_qds_block31_decoder_output	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  divider_1D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_2D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_dffe_1a_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  divider_dffe_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_in_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  padded_2_zeros_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  padded_3_zeros_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  pos_qk0d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk1d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk2d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qkd_mux_input_w :	STD_LOGIC_VECTOR (107 DOWNTO 0);
	 SIGNAL  qkd_mux_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_adder_padded_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_dffe_1a_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  Rk_in_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  Rk_next_dffe_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  rom_add_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  rom_mux_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_1a_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_dffe_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  srt_adder_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int11_w_divider_in_w_range1513w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 COMPONENT  Float_32_Div_altfp_div_csa_lsa
	 PORT
	 ( 
		add_sub	:	IN  STD_LOGIC := '1';
		dataa	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(26 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_qds_block_7o8
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		decoder_bus	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
		decoder_output	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	divider_1D_w <= ( padded_3_zeros_w & "1" & divider_dffe_1a_w);
	divider_2D_w <= ( padded_2_zeros_w & "1" & divider_dffe_1a_w & "0");
	divider_dffe_1a_w <= divider_dffe_1a;
	divider_dffe_w <= ( "1" & divider_dffe);
	divider_in_w <= divider;
	divider_reg <= divider_dffe_w;
	padded_2_zeros_w <= (OTHERS => '0');
	padded_3_zeros_w <= (OTHERS => '0');
	pos_qk0d_int_w <= (OTHERS => '0');
	pos_qk1d_int_w <= divider_1D_w;
	pos_qk2d_int_w <= divider_2D_w;
	qkd_mux_input_w <= ( pos_qk2d_int_w & pos_qk2d_int_w & pos_qk1d_int_w & pos_qk0d_int_w);
	qkd_mux_w <= wire_mux32_result;
	Rk_adder_padded_w <= ( padded_3_zeros_w & Rk_dffe);
	Rk_dffe_1a_w <= Rk_in_w;
	Rk_in_w <= Rk;
	Rk_next <= Rk_next_dffe_w;
	Rk_next_dffe_w <= Rk_next_dffe;
	rom <= rom_out_dffe_w;
	rom_add_w <= ( padded_3_zeros_w & Rk_in_w(23 DOWNTO 19) & divider_in_w(22 DOWNTO 19));
	rom_mux_w <= rom_out_1a_w;
	rom_out_1a_w <= wire_qds_block31_decoder_output;
	rom_out_dffe_w <= rom_out_dffe;
	srt_adder_w <= wire_altfp_div_csa33_result(24 DOWNTO 0);
	wire_srt_block_int11_w_divider_in_w_range1513w <= divider_in_w(22 DOWNTO 0);
	altfp_div_csa33 :  Float_32_Div_altfp_div_csa_lsa
	  PORT MAP ( 
		add_sub => rom_mux_w(2),
		dataa => Rk_adder_padded_w,
		datab => qkd_mux_w,
		result => wire_altfp_div_csa33_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_dffe <= divider_dffe_1a_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_dffe_1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_dffe_1a <= wire_srt_block_int11_w_divider_in_w_range1513w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_dffe <= Rk_dffe_1a_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_next_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_next_dffe <= srt_adder_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_out_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_out_dffe <= rom_out_1a_w;
			END IF;
		END IF;
	END PROCESS;
	loop5 : FOR i IN 0 TO 3 GENERATE
		loop6 : FOR j IN 0 TO 26 GENERATE
			wire_mux32_data_2d(i, j) <= qkd_mux_input_w(i*27+j);
		END GENERATE loop6;
	END GENERATE loop5;
	mux32 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 4,
		LPM_WIDTH => 27,
		LPM_WIDTHS => 2
	  )
	  PORT MAP ( 
		data => wire_mux32_data_2d,
		result => wire_mux32_result,
		sel => rom_mux_w(1 DOWNTO 0)
	  );
	qds_block31 :  Float_32_Div_qds_block_7o8
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		decoder_bus => rom_add_w,
		decoder_output => wire_qds_block31_decoder_output
	  );

 END RTL; --Float_32_Div_srt_block_int_sfk


--srt_block_int CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" OPTIMIZE="AREA" POSITION="MIDDLE" WIDTH_DIV=24 WIDTH_RK_IN=25 WIDTH_RK_OUT=25 WIDTH_ROM=3 WIDTH_ROM_ADD=12 aclr clken clock divider divider_reg Rk Rk_next rom
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END


--qds_block CBX_AUTO_BLACKBOX="ALL" aclr clken clock decoder_bus decoder_output
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_compare 4 lpm_mux 1 reg 3 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_qds_block_6a7 IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 decoder_bus	:	IN  STD_LOGIC_VECTOR (11 DOWNTO 0);
		 decoder_output	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END Float_32_Div_qds_block_6a7;

 ARCHITECTURE RTL OF Float_32_Div_qds_block_6a7 IS

	 SIGNAL	 q_next_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_cmpr44_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr45_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr46_aleb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr47_aleb	:	STD_LOGIC;
	 SIGNAL  wire_mux43_data_2d	:	STD_LOGIC_2D(15 DOWNTO 0, 31 DOWNTO 0);
	 SIGNAL  wire_mux43_result	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_k_comp_w_range1717w1726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_k_comp_w_range1719w1728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_k_comp_w_range1715w1725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_k_comp_w_range1718w1727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_k_comp_w_range1719w1722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1728w1729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1722w1723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  decoder_output_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  Div_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  k_comp_w :	STD_LOGIC_VECTOR (3 DOWNTO 0);
	 SIGNAL  mk_bus_const_w :	STD_LOGIC_VECTOR (511 DOWNTO 0);
	 SIGNAL  mk_bus_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mk_neg1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos0_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  mk_pos2_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  q_next_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  Rk_in_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  Rk_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_k_comp_w_range1715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_k_comp_w_range1717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_k_comp_w_range1718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_qds_block40_w_k_comp_w_range1719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	wire_qds_block40_w_lg_w_k_comp_w_range1717w1726w(0) <= wire_qds_block40_w_k_comp_w_range1717w(0) AND wire_qds_block40_w_lg_w_k_comp_w_range1715w1725w(0);
	wire_qds_block40_w_lg_w_k_comp_w_range1719w1728w(0) <= wire_qds_block40_w_k_comp_w_range1719w(0) AND wire_qds_block40_w_lg_w_k_comp_w_range1718w1727w(0);
	wire_qds_block40_w_lg_w_k_comp_w_range1715w1725w(0) <= NOT wire_qds_block40_w_k_comp_w_range1715w(0);
	wire_qds_block40_w_lg_w_k_comp_w_range1718w1727w(0) <= NOT wire_qds_block40_w_k_comp_w_range1718w(0);
	wire_qds_block40_w_lg_w_k_comp_w_range1719w1722w(0) <= NOT wire_qds_block40_w_k_comp_w_range1719w(0);
	wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1728w1729w(0) <= wire_qds_block40_w_lg_w_k_comp_w_range1719w1728w(0) OR wire_qds_block40_w_lg_w_k_comp_w_range1717w1726w(0);
	wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1722w1723w(0) <= wire_qds_block40_w_lg_w_k_comp_w_range1719w1722w(0) OR wire_qds_block40_w_k_comp_w_range1715w(0);
	decoder_output <= decoder_output_w;
	decoder_output_w <= q_next_dffe;
	Div_w <= decoder_bus(3 DOWNTO 0);
	k_comp_w <= ( wire_cmpr47_aleb & wire_cmpr46_aleb & wire_cmpr45_aleb & wire_cmpr44_aleb);
	mk_bus_const_w <= ( "01011101000111111110000110100011" & "01011010000111101110001010100110" & "01010111000111011110001110101001" & "01010100000111001110010010101100" & "01010001000110111110010110101111" & "01001110000110101110011010110010" & "01001011000110011110011110110101" & "01001000000110001110100010111000" & "01000101000101111110100110111011" & "01000010000101101110101010111110" & "00111111000101011110101111000001" & "00111100000101001110110011000100" & "00111001000100111110110111000111" & "00110110000100101110111011001010" & "00110011000100011110111111001101" & "00110000000100001111000011010000");
	mk_bus_w <= wire_mux43_result;
	mk_neg1_w <= ( mk_bus_w(7) & mk_bus_w(7 DOWNTO 0));
	mk_pos0_w <= ( mk_bus_w(15) & mk_bus_w(15 DOWNTO 8));
	mk_pos1_w <= ( mk_bus_w(23) & mk_bus_w(23 DOWNTO 16));
	mk_pos2_w <= ( mk_bus_w(31) & mk_bus_w(31 DOWNTO 24));
	q_next_w <= ( k_comp_w(1) & wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1722w1723w & wire_qds_block40_w_lg_w_lg_w_k_comp_w_range1719w1728w1729w);
	Rk_in_w <= ( decoder_bus(11 DOWNTO 4) & "0");
	Rk_w <= Rk_in_w;
	wire_qds_block40_w_k_comp_w_range1715w(0) <= k_comp_w(0);
	wire_qds_block40_w_k_comp_w_range1717w(0) <= k_comp_w(1);
	wire_qds_block40_w_k_comp_w_range1718w(0) <= k_comp_w(2);
	wire_qds_block40_w_k_comp_w_range1719w(0) <= k_comp_w(3);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN q_next_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN q_next_dffe <= q_next_w;
			END IF;
		END IF;
	END PROCESS;
	cmpr44 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr44_aleb,
		dataa => Rk_w,
		datab => mk_neg1_w
	  );
	cmpr45 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr45_aleb,
		dataa => Rk_w,
		datab => mk_pos0_w
	  );
	cmpr46 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr46_aleb,
		dataa => Rk_w,
		datab => mk_pos1_w
	  );
	cmpr47 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aleb => wire_cmpr47_aleb,
		dataa => Rk_w,
		datab => mk_pos2_w
	  );
	loop7 : FOR i IN 0 TO 15 GENERATE
		loop8 : FOR j IN 0 TO 31 GENERATE
			wire_mux43_data_2d(i, j) <= mk_bus_const_w(i*32+j);
		END GENERATE loop8;
	END GENERATE loop7;
	mux43 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 16,
		LPM_WIDTH => 32,
		LPM_WIDTHS => 4
	  )
	  PORT MAP ( 
		data => wire_mux43_data_2d,
		result => wire_mux43_result,
		sel => Div_w
	  );

 END RTL; --Float_32_Div_qds_block_6a7

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 1 lpm_compare 4 lpm_mux 2 reg 102 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_srt_block_int_4ik IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 divider	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 divider_reg	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 Rk	:	IN  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 Rk_next	:	OUT  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 rom	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END Float_32_Div_srt_block_int_4ik;

 ARCHITECTURE RTL OF Float_32_Div_srt_block_int_4ik IS

	 SIGNAL  wire_altfp_div_csa42_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL	 divider_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 divider_dffe_1a	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_dffe	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_next_dffe	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_out_dffe	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mux41_data_2d	:	STD_LOGIC_2D(3 DOWNTO 0, 26 DOWNTO 0);
	 SIGNAL  wire_mux41_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_qds_block40_decoder_output	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  divider_1D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_2D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_dffe_1a_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  divider_dffe_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_in_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  padded_2_zeros_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  padded_3_zeros_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  pos_qk0d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk1d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk2d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qkd_mux_input_w :	STD_LOGIC_VECTOR (107 DOWNTO 0);
	 SIGNAL  qkd_mux_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_adder_padded_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_dffe_1a_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_in_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_dffe_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  rom_add_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  rom_mux_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_1a_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_dffe_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  srt_adder_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int12_w_divider_in_w_range1628w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 COMPONENT  Float_32_Div_altfp_div_csa_lsa
	 PORT
	 ( 
		add_sub	:	IN  STD_LOGIC := '1';
		dataa	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(26 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_qds_block_6a7
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		decoder_bus	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
		decoder_output	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	divider_1D_w <= ( padded_3_zeros_w & "1" & divider_dffe_1a_w);
	divider_2D_w <= ( padded_2_zeros_w & "1" & divider_dffe_1a_w & "0");
	divider_dffe_1a_w <= divider_dffe_1a;
	divider_dffe_w <= ( "1" & divider_dffe);
	divider_in_w <= divider;
	divider_reg <= divider_dffe_w;
	padded_2_zeros_w <= (OTHERS => '0');
	padded_3_zeros_w <= (OTHERS => '0');
	pos_qk0d_int_w <= (OTHERS => '0');
	pos_qk1d_int_w <= divider_1D_w;
	pos_qk2d_int_w <= divider_2D_w;
	qkd_mux_input_w <= ( pos_qk2d_int_w & pos_qk2d_int_w & pos_qk1d_int_w & pos_qk0d_int_w);
	qkd_mux_w <= wire_mux41_result;
	Rk_adder_padded_w <= ( Rk_dffe & padded_2_zeros_w);
	Rk_dffe_1a_w <= Rk_in_w;
	Rk_in_w <= Rk;
	Rk_next <= Rk_next_dffe_w;
	Rk_next_dffe_w <= Rk_next_dffe;
	rom <= rom_out_dffe_w;
	rom_add_w <= ( Rk_in_w(24 DOWNTO 17) & divider_in_w(22 DOWNTO 19));
	rom_mux_w <= rom_out_1a_w;
	rom_out_1a_w <= wire_qds_block40_decoder_output;
	rom_out_dffe_w <= rom_out_dffe;
	srt_adder_w <= wire_altfp_div_csa42_result(24 DOWNTO 0);
	wire_srt_block_int12_w_divider_in_w_range1628w <= divider_in_w(22 DOWNTO 0);
	altfp_div_csa42 :  Float_32_Div_altfp_div_csa_lsa
	  PORT MAP ( 
		add_sub => rom_mux_w(2),
		dataa => Rk_adder_padded_w,
		datab => qkd_mux_w,
		result => wire_altfp_div_csa42_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_dffe <= divider_dffe_1a_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_dffe_1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_dffe_1a <= wire_srt_block_int12_w_divider_in_w_range1628w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_dffe <= Rk_dffe_1a_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_next_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_next_dffe <= srt_adder_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_out_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_out_dffe <= rom_out_1a_w;
			END IF;
		END IF;
	END PROCESS;
	loop9 : FOR i IN 0 TO 3 GENERATE
		loop10 : FOR j IN 0 TO 26 GENERATE
			wire_mux41_data_2d(i, j) <= qkd_mux_input_w(i*27+j);
		END GENERATE loop10;
	END GENERATE loop9;
	mux41 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 4,
		LPM_WIDTH => 27,
		LPM_WIDTHS => 2
	  )
	  PORT MAP ( 
		data => wire_mux41_data_2d,
		result => wire_mux41_result,
		sel => rom_mux_w(1 DOWNTO 0)
	  );
	qds_block40 :  Float_32_Div_qds_block_6a7
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		decoder_bus => rom_add_w,
		decoder_output => wire_qds_block40_decoder_output
	  );

 END RTL; --Float_32_Div_srt_block_int_4ik


--srt_block_int CBX_AUTO_BLACKBOX="ALL" DEVICE_FAMILY="Cyclone IV E" OPTIMIZE="AREA" POSITION="LAST" WIDTH_DIV=24 WIDTH_RK_IN=25 WIDTH_RK_OUT=27 WIDTH_ROM=3 WIDTH_ROM_ADD=12 aclr clken clock divider divider_reg Rk Rk_next rom
--VERSION_BEGIN 18.1 cbx_altbarrel_shift 2018:09:12:13:04:09:SJ cbx_altera_syncram_nd_impl 2018:09:12:13:04:09:SJ cbx_altfp_div 2018:09:12:13:04:09:SJ cbx_altsyncram 2018:09:12:13:04:09:SJ cbx_cycloneii 2018:09:12:13:04:09:SJ cbx_lpm_abs 2018:09:12:13:04:09:SJ cbx_lpm_add_sub 2018:09:12:13:04:09:SJ cbx_lpm_compare 2018:09:12:13:04:09:SJ cbx_lpm_decode 2018:09:12:13:04:09:SJ cbx_lpm_divide 2018:09:12:13:04:09:SJ cbx_lpm_mult 2018:09:12:13:04:09:SJ cbx_lpm_mux 2018:09:12:13:04:09:SJ cbx_mgl 2018:09:12:14:15:07:SJ cbx_nadder 2018:09:12:13:04:09:SJ cbx_padd 2018:09:12:13:04:09:SJ cbx_stratix 2018:09:12:13:04:09:SJ cbx_stratixii 2018:09:12:13:04:09:SJ cbx_stratixiii 2018:09:12:13:04:09:SJ cbx_stratixv 2018:09:12:13:04:09:SJ cbx_util_mgl 2018:09:12:13:04:09:SJ  VERSION_END

 LIBRARY lpm;
 USE lpm.lpm_components.all;

--synthesis_resources = lpm_add_sub 1 lpm_compare 4 lpm_mux 2 reg 51 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_srt_block_int_bck IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 divider	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 divider_reg	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 Rk	:	IN  STD_LOGIC_VECTOR (24 DOWNTO 0);
		 Rk_next	:	OUT  STD_LOGIC_VECTOR (26 DOWNTO 0);
		 rom	:	OUT  STD_LOGIC_VECTOR (2 DOWNTO 0)
	 ); 
 END Float_32_Div_srt_block_int_bck;

 ARCHITECTURE RTL OF Float_32_Div_srt_block_int_bck IS

	 SIGNAL  wire_altfp_div_csa50_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL	 divider_dffe_1a	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_dffe	:	STD_LOGIC_VECTOR(24 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_mux49_data_2d	:	STD_LOGIC_2D(3 DOWNTO 0, 26 DOWNTO 0);
	 SIGNAL  wire_mux49_result	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_qds_block48_decoder_output	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  divider_1D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_2D_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  divider_dffe_1a_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  divider_dffe_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_in_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  padded_2_zeros_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  padded_3_zeros_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  pos_qk0d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk1d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  pos_qk2d_int_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  qkd_mux_input_w :	STD_LOGIC_VECTOR (107 DOWNTO 0);
	 SIGNAL  qkd_mux_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_adder_padded_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_dffe_1a_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_in_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_dffe_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  rom_add_w :	STD_LOGIC_VECTOR (11 DOWNTO 0);
	 SIGNAL  rom_mux_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_1a_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_dffe_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  srt_adder_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_srt_block_int24_w_divider_in_w_range1738w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 COMPONENT  Float_32_Div_altfp_div_csa_lsa
	 PORT
	 ( 
		add_sub	:	IN  STD_LOGIC := '1';
		dataa	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(26 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(26 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_qds_block_6a7
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		decoder_bus	:	IN  STD_LOGIC_VECTOR(11 DOWNTO 0);
		decoder_output	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	divider_1D_w <= ( padded_3_zeros_w & "1" & divider_dffe_1a_w);
	divider_2D_w <= ( padded_2_zeros_w & "1" & divider_dffe_1a_w & "0");
	divider_dffe_1a_w <= divider_dffe_1a;
	divider_dffe_w <= ( "1" & divider_dffe_1a_w);
	divider_in_w <= divider;
	divider_reg <= divider_dffe_w;
	padded_2_zeros_w <= (OTHERS => '0');
	padded_3_zeros_w <= (OTHERS => '0');
	pos_qk0d_int_w <= (OTHERS => '0');
	pos_qk1d_int_w <= divider_1D_w;
	pos_qk2d_int_w <= divider_2D_w;
	qkd_mux_input_w <= ( pos_qk2d_int_w & pos_qk2d_int_w & pos_qk1d_int_w & pos_qk0d_int_w);
	qkd_mux_w <= wire_mux49_result;
	Rk_adder_padded_w <= ( Rk_dffe & padded_2_zeros_w);
	Rk_dffe_1a_w <= Rk_in_w;
	Rk_in_w <= Rk;
	Rk_next <= Rk_next_dffe_w;
	Rk_next_dffe_w <= srt_adder_w;
	rom <= rom_out_dffe_w;
	rom_add_w <= ( Rk_in_w(24 DOWNTO 17) & divider_in_w(22 DOWNTO 19));
	rom_mux_w <= rom_out_1a_w;
	rom_out_1a_w <= wire_qds_block48_decoder_output;
	rom_out_dffe_w <= rom_out_1a_w;
	srt_adder_w <= wire_altfp_div_csa50_result(26 DOWNTO 0);
	wire_srt_block_int24_w_divider_in_w_range1738w <= divider_in_w(22 DOWNTO 0);
	altfp_div_csa50 :  Float_32_Div_altfp_div_csa_lsa
	  PORT MAP ( 
		add_sub => rom_mux_w(2),
		dataa => Rk_adder_padded_w,
		datab => qkd_mux_w,
		result => wire_altfp_div_csa50_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_dffe_1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_dffe_1a <= wire_srt_block_int24_w_divider_in_w_range1738w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_dffe <= Rk_dffe_1a_w;
			END IF;
		END IF;
	END PROCESS;
	loop11 : FOR i IN 0 TO 3 GENERATE
		loop12 : FOR j IN 0 TO 26 GENERATE
			wire_mux49_data_2d(i, j) <= qkd_mux_input_w(i*27+j);
		END GENERATE loop12;
	END GENERATE loop11;
	mux49 :  lpm_mux
	  GENERIC MAP (
		LPM_SIZE => 4,
		LPM_WIDTH => 27,
		LPM_WIDTHS => 2
	  )
	  PORT MAP ( 
		data => wire_mux49_data_2d,
		result => wire_mux49_result,
		sel => rom_mux_w(1 DOWNTO 0)
	  );
	qds_block48 :  Float_32_Div_qds_block_6a7
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		decoder_bus => rom_add_w,
		decoder_output => wire_qds_block48_decoder_output
	  );

 END RTL; --Float_32_Div_srt_block_int_bck

--synthesis_resources = lpm_add_sub 17 lpm_compare 56 lpm_mux 28 reg 1908 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_srt_ext_14f IS 
	 PORT 
	 ( 
		 aclr	:	IN  STD_LOGIC := '0';
		 clken	:	IN  STD_LOGIC := '1';
		 clock	:	IN  STD_LOGIC := '0';
		 denom	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 divider	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 numer	:	IN  STD_LOGIC_VECTOR (23 DOWNTO 0);
		 quotient	:	OUT  STD_LOGIC_VECTOR (27 DOWNTO 0);
		 remain	:	OUT  STD_LOGIC_VECTOR (23 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_srt_ext_14f;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_srt_ext_14f IS

	 SIGNAL  wire_altfp_div_csa25_result	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_csa26_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altfp_div_csa27_result	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL	 divider_next_special_dffe	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 Rk_remainder_special_dffe	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe0c	:	STD_LOGIC_VECTOR(49 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe10c	:	STD_LOGIC_VECTOR(14 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe11c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe12c	:	STD_LOGIC_VECTOR(2 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe1c	:	STD_LOGIC_VECTOR(68 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe2c	:	STD_LOGIC_VECTOR(62 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe3c	:	STD_LOGIC_VECTOR(56 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe4c	:	STD_LOGIC_VECTOR(50 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe5c	:	STD_LOGIC_VECTOR(44 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe6c	:	STD_LOGIC_VECTOR(38 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe7c	:	STD_LOGIC_VECTOR(32 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe8c	:	STD_LOGIC_VECTOR(26 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rom_reg_dffe9c	:	STD_LOGIC_VECTOR(20 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_srt_block_int11_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int11_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int11_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int12_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int12_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int12_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int13_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int13_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int13_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int14_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int14_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int14_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int15_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int15_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int15_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int16_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int16_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int16_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int17_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int17_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int17_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int18_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int18_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int18_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int19_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int19_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int19_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int20_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int20_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int20_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int21_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int21_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int21_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int22_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int22_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int22_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int23_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int23_Rk_next	:	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  wire_srt_block_int23_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_srt_block_int24_divider_reg	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_srt_block_int24_Rk_next	:	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  wire_srt_block_int24_rom	:	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1504w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1501w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1422w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1353w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1452w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1403w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1455w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1408w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1458w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1413w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1461w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1418w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1425w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1358w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1428w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1363w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1431w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1368w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1434w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1373w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1437w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1378w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1440w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1383w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1443w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1388w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1446w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1393w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1449w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1398w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1499w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1503w	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1354w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1421w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1404w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1451w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1409w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1454w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1414w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1457w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1419w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1460w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1359w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1424w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1364w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1427w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1369w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1430w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1374w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1433w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1379w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1436w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1384w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1439w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1389w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1442w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1394w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1445w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1399w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1448w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1352w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1402w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1407w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1417w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1357w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1362w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1367w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1372w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1377w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1382w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1387w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1392w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1397w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  added_remainder_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_dffe_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_special_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w0c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w10c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w11c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w12c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w13c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w1c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w2c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w3c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w4c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w5c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w6c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w7c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w8c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_next_w9c :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  divider_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  full_neg_rom_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  full_pos_rom_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  mux_remainder_w :	STD_LOGIC;
	 SIGNAL  neg_rom_w0c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w10c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w11c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w12c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w13c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w1c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w2c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w3c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w4c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w5c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w6c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w7c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w8c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  neg_rom_w9c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w0c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w10c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w11c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w12c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w13c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w1c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w2c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w3c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w4c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w5c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w6c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w7c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w8c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  pos_rom_w9c :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  Rk_next0_w :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w0c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w10c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w11c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w12c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w13c :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_next_w1c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w2c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w3c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w4c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w5c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w6c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w7c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w8c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_next_w9c :	STD_LOGIC_VECTOR (24 DOWNTO 0);
	 SIGNAL  Rk_remainder_special_w :	STD_LOGIC_VECTOR (26 DOWNTO 0);
	 SIGNAL  Rk_remainder_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  Rk_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  rom_dffe_w0c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w10c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w11c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w12c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w13c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w1c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w2c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w3c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w4c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w5c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w6c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w7c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w8c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_dffe_w9c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_mux_w :	STD_LOGIC_VECTOR (13 DOWNTO 0);
	 SIGNAL  rom_out_1a_w :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w0c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w10c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w11c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w12c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w13c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w1c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w2c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w3c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w4c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w5c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w6c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w7c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w8c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  rom_out_w9c :	STD_LOGIC_VECTOR (2 DOWNTO 0);
	 SIGNAL  srt_adjust_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  srt_adjusted_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  true_quotient_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  value_one_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  zero_quotient_w :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_Rk_remainder_special_w_range1498w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w0c_range1311w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w10c_range1401w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w11c_range1406w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w12c_range1411w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w13c_range1416w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w1c_range1356w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w2c_range1361w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w3c_range1366w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w4c_range1371w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w5c_range1376w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w6c_range1381w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w7c_range1386w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w8c_range1391w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_dffe_w9c_range1396w	:	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1324w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1349w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1351w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1331w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1341w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_w_rom_mux_w_range1343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  Float_32_Div_altfp_div_csa_jub
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_altfp_div_csa_vse
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		dataa	:	IN  STD_LOGIC_VECTOR(27 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(27 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(27 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_altfp_div_csa_ovb
	 PORT
	 ( 
		dataa	:	IN  STD_LOGIC_VECTOR(27 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(27 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(27 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_srt_block_int_sfk
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		divider	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		divider_reg	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0);
		Rk	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		Rk_next	:	OUT  STD_LOGIC_VECTOR(24 DOWNTO 0);
		rom	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_srt_block_int_4ik
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		divider	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		divider_reg	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0);
		Rk	:	IN  STD_LOGIC_VECTOR(24 DOWNTO 0);
		Rk_next	:	OUT  STD_LOGIC_VECTOR(24 DOWNTO 0);
		rom	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_srt_block_int_bck
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		divider	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		divider_reg	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0);
		Rk	:	IN  STD_LOGIC_VECTOR(24 DOWNTO 0);
		Rk_next	:	OUT  STD_LOGIC_VECTOR(26 DOWNTO 0);
		rom	:	OUT  STD_LOGIC_VECTOR(2 DOWNTO 0)
	 ); 
	 END COMPONENT;
 BEGIN

	loop13 : FOR i IN 0 TO 27 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1504w(i) <= wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1500w(0) AND srt_adjust_w(i);
	END GENERATE loop13;
	loop14 : FOR i IN 0 TO 23 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1501w(i) <= wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1500w(0) AND wire_altfp_div_srt_ext1_w_Rk_remainder_special_w_range1498w(i);
	END GENERATE loop14;
	loop15 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1422w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1352w(0) AND zero_quotient_w(i);
	END GENERATE loop15;
	loop16 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1353w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1352w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w0c_range1311w(i);
	END GENERATE loop16;
	loop17 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1452w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1402w(0) AND zero_quotient_w(i);
	END GENERATE loop17;
	loop18 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1403w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1402w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w10c_range1401w(i);
	END GENERATE loop18;
	loop19 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1455w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1407w(0) AND zero_quotient_w(i);
	END GENERATE loop19;
	loop20 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1408w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1407w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w11c_range1406w(i);
	END GENERATE loop20;
	loop21 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1458w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1412w(0) AND zero_quotient_w(i);
	END GENERATE loop21;
	loop22 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1413w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1412w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w12c_range1411w(i);
	END GENERATE loop22;
	loop23 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1461w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1417w(0) AND zero_quotient_w(i);
	END GENERATE loop23;
	loop24 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1418w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1417w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w13c_range1416w(i);
	END GENERATE loop24;
	loop25 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1425w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1357w(0) AND zero_quotient_w(i);
	END GENERATE loop25;
	loop26 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1358w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1357w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w1c_range1356w(i);
	END GENERATE loop26;
	loop27 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1428w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1362w(0) AND zero_quotient_w(i);
	END GENERATE loop27;
	loop28 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1363w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1362w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w2c_range1361w(i);
	END GENERATE loop28;
	loop29 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1431w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1367w(0) AND zero_quotient_w(i);
	END GENERATE loop29;
	loop30 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1368w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1367w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w3c_range1366w(i);
	END GENERATE loop30;
	loop31 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1434w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1372w(0) AND zero_quotient_w(i);
	END GENERATE loop31;
	loop32 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1373w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1372w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w4c_range1371w(i);
	END GENERATE loop32;
	loop33 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1437w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1377w(0) AND zero_quotient_w(i);
	END GENERATE loop33;
	loop34 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1378w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1377w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w5c_range1376w(i);
	END GENERATE loop34;
	loop35 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1440w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1382w(0) AND zero_quotient_w(i);
	END GENERATE loop35;
	loop36 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1383w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1382w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w6c_range1381w(i);
	END GENERATE loop36;
	loop37 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1443w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1387w(0) AND zero_quotient_w(i);
	END GENERATE loop37;
	loop38 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1388w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1387w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w7c_range1386w(i);
	END GENERATE loop38;
	loop39 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1446w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1392w(0) AND zero_quotient_w(i);
	END GENERATE loop39;
	loop40 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1393w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1392w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w8c_range1391w(i);
	END GENERATE loop40;
	loop41 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1449w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1397w(0) AND zero_quotient_w(i);
	END GENERATE loop41;
	loop42 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1398w(i) <= wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1397w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w9c_range1396w(i);
	END GENERATE loop42;
	loop43 : FOR i IN 0 TO 23 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1499w(i) <= mux_remainder_w AND added_remainder_w(i);
	END GENERATE loop43;
	loop44 : FOR i IN 0 TO 27 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1503w(i) <= mux_remainder_w AND srt_adjusted_w(i);
	END GENERATE loop44;
	loop45 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1354w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1324w(0) AND zero_quotient_w(i);
	END GENERATE loop45;
	loop46 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1421w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1324w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w0c_range1311w(i);
	END GENERATE loop46;
	loop47 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1404w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1345w(0) AND zero_quotient_w(i);
	END GENERATE loop47;
	loop48 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1451w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1345w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w10c_range1401w(i);
	END GENERATE loop48;
	loop49 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1409w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1347w(0) AND zero_quotient_w(i);
	END GENERATE loop49;
	loop50 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1454w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1347w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w11c_range1406w(i);
	END GENERATE loop50;
	loop51 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1414w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1349w(0) AND zero_quotient_w(i);
	END GENERATE loop51;
	loop52 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1457w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1349w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w12c_range1411w(i);
	END GENERATE loop52;
	loop53 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1419w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1351w(0) AND zero_quotient_w(i);
	END GENERATE loop53;
	loop54 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1460w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1351w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w13c_range1416w(i);
	END GENERATE loop54;
	loop55 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1359w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1327w(0) AND zero_quotient_w(i);
	END GENERATE loop55;
	loop56 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1424w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1327w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w1c_range1356w(i);
	END GENERATE loop56;
	loop57 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1364w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1329w(0) AND zero_quotient_w(i);
	END GENERATE loop57;
	loop58 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1427w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1329w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w2c_range1361w(i);
	END GENERATE loop58;
	loop59 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1369w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1331w(0) AND zero_quotient_w(i);
	END GENERATE loop59;
	loop60 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1430w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1331w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w3c_range1366w(i);
	END GENERATE loop60;
	loop61 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1374w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1333w(0) AND zero_quotient_w(i);
	END GENERATE loop61;
	loop62 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1433w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1333w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w4c_range1371w(i);
	END GENERATE loop62;
	loop63 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1379w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1335w(0) AND zero_quotient_w(i);
	END GENERATE loop63;
	loop64 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1436w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1335w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w5c_range1376w(i);
	END GENERATE loop64;
	loop65 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1384w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1337w(0) AND zero_quotient_w(i);
	END GENERATE loop65;
	loop66 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1439w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1337w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w6c_range1381w(i);
	END GENERATE loop66;
	loop67 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1389w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1339w(0) AND zero_quotient_w(i);
	END GENERATE loop67;
	loop68 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1442w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1339w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w7c_range1386w(i);
	END GENERATE loop68;
	loop69 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1394w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1341w(0) AND zero_quotient_w(i);
	END GENERATE loop69;
	loop70 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1445w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1341w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w8c_range1391w(i);
	END GENERATE loop70;
	loop71 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1399w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1343w(0) AND zero_quotient_w(i);
	END GENERATE loop71;
	loop72 : FOR i IN 0 TO 1 GENERATE 
		wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1448w(i) <= wire_altfp_div_srt_ext1_w_rom_mux_w_range1343w(0) AND wire_altfp_div_srt_ext1_w_rom_dffe_w9c_range1396w(i);
	END GENERATE loop72;
	wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1500w(0) <= NOT mux_remainder_w;
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1352w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1324w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1402w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1345w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1407w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1347w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1412w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1349w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1417w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1351w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1357w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1327w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1362w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1329w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1367w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1331w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1372w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1333w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1377w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1335w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1382w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1337w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1387w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1339w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1392w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1341w(0);
	wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1397w(0) <= NOT wire_altfp_div_srt_ext1_w_rom_mux_w_range1343w(0);
	added_remainder_w <= wire_altfp_div_csa25_result;
	divider <= divider_next_special_w;
	divider_dffe_w <= wire_srt_block_int11_divider_reg;
	divider_next_special_w <= divider_next_special_dffe;
	divider_next_w0c <= divider_dffe_w;
	divider_next_w10c <= wire_srt_block_int21_divider_reg;
	divider_next_w11c <= wire_srt_block_int22_divider_reg;
	divider_next_w12c <= wire_srt_block_int23_divider_reg;
	divider_next_w13c <= wire_srt_block_int24_divider_reg;
	divider_next_w1c <= wire_srt_block_int12_divider_reg;
	divider_next_w2c <= wire_srt_block_int13_divider_reg;
	divider_next_w3c <= wire_srt_block_int14_divider_reg;
	divider_next_w4c <= wire_srt_block_int15_divider_reg;
	divider_next_w5c <= wire_srt_block_int16_divider_reg;
	divider_next_w6c <= wire_srt_block_int17_divider_reg;
	divider_next_w7c <= wire_srt_block_int18_divider_reg;
	divider_next_w8c <= wire_srt_block_int19_divider_reg;
	divider_next_w9c <= wire_srt_block_int20_divider_reg;
	divider_w <= denom;
	full_neg_rom_w <= ( neg_rom_w0c & neg_rom_w1c & neg_rom_w2c & neg_rom_w3c & neg_rom_w4c & neg_rom_w5c & neg_rom_w6c & neg_rom_w7c & neg_rom_w8c & neg_rom_w9c & neg_rom_w10c & neg_rom_w11c & neg_rom_w12c & neg_rom_w13c);
	full_pos_rom_w <= ( pos_rom_w0c & pos_rom_w1c & pos_rom_w2c & pos_rom_w3c & pos_rom_w4c & pos_rom_w5c & pos_rom_w6c & pos_rom_w7c & pos_rom_w8c & pos_rom_w9c & pos_rom_w10c & pos_rom_w11c & pos_rom_w12c & pos_rom_w13c);
	mux_remainder_w <= ((Rk_remainder_special_w(26) OR Rk_remainder_special_w(25)) OR Rk_remainder_special_w(24));
	neg_rom_w0c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1422w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1421w);
	neg_rom_w10c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1452w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1451w);
	neg_rom_w11c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1455w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1454w);
	neg_rom_w12c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1458w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1457w);
	neg_rom_w13c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1461w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1460w);
	neg_rom_w1c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1425w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1424w);
	neg_rom_w2c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1428w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1427w);
	neg_rom_w3c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1431w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1430w);
	neg_rom_w4c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1434w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1433w);
	neg_rom_w5c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1437w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1436w);
	neg_rom_w6c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1440w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1439w);
	neg_rom_w7c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1443w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1442w);
	neg_rom_w8c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1446w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1445w);
	neg_rom_w9c <= (wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1449w OR wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1448w);
	pos_rom_w0c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1324w1354w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1324w1352w1353w);
	pos_rom_w10c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1345w1404w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1345w1402w1403w);
	pos_rom_w11c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1347w1409w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1347w1407w1408w);
	pos_rom_w12c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1349w1414w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1349w1412w1413w);
	pos_rom_w13c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1351w1419w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1351w1417w1418w);
	pos_rom_w1c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1327w1359w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1327w1357w1358w);
	pos_rom_w2c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1329w1364w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1329w1362w1363w);
	pos_rom_w3c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1331w1369w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1331w1367w1368w);
	pos_rom_w4c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1333w1374w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1333w1372w1373w);
	pos_rom_w5c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1335w1379w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1335w1377w1378w);
	pos_rom_w6c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1337w1384w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1337w1382w1383w);
	pos_rom_w7c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1339w1389w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1339w1387w1388w);
	pos_rom_w8c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1341w1394w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1341w1392w1393w);
	pos_rom_w9c <= (wire_altfp_div_srt_ext1_w_lg_w_rom_mux_w_range1343w1399w OR wire_altfp_div_srt_ext1_w_lg_w_lg_w_rom_mux_w_range1343w1397w1398w);
	quotient <= true_quotient_w;
	remain <= Rk_remainder_w;
	Rk_next0_w <= wire_srt_block_int11_Rk_next;
	Rk_next_w0c <= Rk_next0_w;
	Rk_next_w10c <= wire_srt_block_int21_Rk_next;
	Rk_next_w11c <= wire_srt_block_int22_Rk_next;
	Rk_next_w12c <= wire_srt_block_int23_Rk_next;
	Rk_next_w13c <= wire_srt_block_int24_Rk_next;
	Rk_next_w1c <= wire_srt_block_int12_Rk_next;
	Rk_next_w2c <= wire_srt_block_int13_Rk_next;
	Rk_next_w3c <= wire_srt_block_int14_Rk_next;
	Rk_next_w4c <= wire_srt_block_int15_Rk_next;
	Rk_next_w5c <= wire_srt_block_int16_Rk_next;
	Rk_next_w6c <= wire_srt_block_int17_Rk_next;
	Rk_next_w7c <= wire_srt_block_int18_Rk_next;
	Rk_next_w8c <= wire_srt_block_int19_Rk_next;
	Rk_next_w9c <= wire_srt_block_int20_Rk_next;
	Rk_remainder_special_w <= Rk_remainder_special_dffe;
	Rk_remainder_w <= (wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1501w OR wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1499w);
	Rk_w <= numer;
	rom_dffe_w0c <= ( "0" & rom_reg_dffe0c(49 DOWNTO 48));
	rom_dffe_w10c <= rom_reg_dffe10c(14 DOWNTO 12);
	rom_dffe_w11c <= rom_reg_dffe11c(8 DOWNTO 6);
	rom_dffe_w12c <= rom_reg_dffe12c(2 DOWNTO 0);
	rom_dffe_w13c <= rom_out_w13c;
	rom_dffe_w1c <= rom_reg_dffe1c(68 DOWNTO 66);
	rom_dffe_w2c <= rom_reg_dffe2c(62 DOWNTO 60);
	rom_dffe_w3c <= rom_reg_dffe3c(56 DOWNTO 54);
	rom_dffe_w4c <= rom_reg_dffe4c(50 DOWNTO 48);
	rom_dffe_w5c <= rom_reg_dffe5c(44 DOWNTO 42);
	rom_dffe_w6c <= rom_reg_dffe6c(38 DOWNTO 36);
	rom_dffe_w7c <= rom_reg_dffe7c(32 DOWNTO 30);
	rom_dffe_w8c <= rom_reg_dffe8c(26 DOWNTO 24);
	rom_dffe_w9c <= rom_reg_dffe9c(20 DOWNTO 18);
	rom_mux_w <= ( rom_dffe_w13c(2) & rom_dffe_w12c(2) & rom_dffe_w11c(2) & rom_dffe_w10c(2) & rom_dffe_w9c(2) & rom_dffe_w8c(2) & rom_dffe_w7c(2) & rom_dffe_w6c(2) & rom_dffe_w5c(2) & rom_dffe_w4c(2) & rom_dffe_w3c(2) & rom_dffe_w2c(2) & rom_dffe_w1c(2) & rom_dffe_w0c(2));
	rom_out_1a_w <= wire_srt_block_int11_rom;
	rom_out_w0c <= rom_out_1a_w;
	rom_out_w10c <= wire_srt_block_int21_rom;
	rom_out_w11c <= wire_srt_block_int22_rom;
	rom_out_w12c <= wire_srt_block_int23_rom;
	rom_out_w13c <= wire_srt_block_int24_rom;
	rom_out_w1c <= wire_srt_block_int12_rom;
	rom_out_w2c <= wire_srt_block_int13_rom;
	rom_out_w3c <= wire_srt_block_int14_rom;
	rom_out_w4c <= wire_srt_block_int15_rom;
	rom_out_w5c <= wire_srt_block_int16_rom;
	rom_out_w6c <= wire_srt_block_int17_rom;
	rom_out_w7c <= wire_srt_block_int18_rom;
	rom_out_w8c <= wire_srt_block_int19_rom;
	rom_out_w9c <= wire_srt_block_int20_rom;
	srt_adjust_w <= wire_altfp_div_csa26_result;
	srt_adjusted_w <= wire_altfp_div_csa27_result;
	true_quotient_w <= (wire_altfp_div_srt_ext1_w_lg_w_lg_mux_remainder_w1500w1504w OR wire_altfp_div_srt_ext1_w_lg_mux_remainder_w1503w);
	value_one_w <= "0000000000000000000000000001";
	zero_quotient_w <= (OTHERS => '0');
	wire_altfp_div_srt_ext1_w_Rk_remainder_special_w_range1498w <= Rk_remainder_special_w(23 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w0c_range1311w <= rom_dffe_w0c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w10c_range1401w <= rom_dffe_w10c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w11c_range1406w <= rom_dffe_w11c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w12c_range1411w <= rom_dffe_w12c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w13c_range1416w <= rom_dffe_w13c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w1c_range1356w <= rom_dffe_w1c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w2c_range1361w <= rom_dffe_w2c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w3c_range1366w <= rom_dffe_w3c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w4c_range1371w <= rom_dffe_w4c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w5c_range1376w <= rom_dffe_w5c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w6c_range1381w <= rom_dffe_w6c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w7c_range1386w <= rom_dffe_w7c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w8c_range1391w <= rom_dffe_w8c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_dffe_w9c_range1396w <= rom_dffe_w9c(1 DOWNTO 0);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1324w(0) <= rom_mux_w(0);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1345w(0) <= rom_mux_w(10);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1347w(0) <= rom_mux_w(11);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1349w(0) <= rom_mux_w(12);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1351w(0) <= rom_mux_w(13);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1327w(0) <= rom_mux_w(1);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1329w(0) <= rom_mux_w(2);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1331w(0) <= rom_mux_w(3);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1333w(0) <= rom_mux_w(4);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1335w(0) <= rom_mux_w(5);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1337w(0) <= rom_mux_w(6);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1339w(0) <= rom_mux_w(7);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1341w(0) <= rom_mux_w(8);
	wire_altfp_div_srt_ext1_w_rom_mux_w_range1343w(0) <= rom_mux_w(9);
	altfp_div_csa25 :  Float_32_Div_altfp_div_csa_jub
	  PORT MAP ( 
		dataa => Rk_remainder_special_w(23 DOWNTO 0),
		datab => divider_next_special_w,
		result => wire_altfp_div_csa25_result
	  );
	altfp_div_csa26 :  Float_32_Div_altfp_div_csa_vse
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		dataa => full_pos_rom_w,
		datab => full_neg_rom_w,
		result => wire_altfp_div_csa26_result
	  );
	altfp_div_csa27 :  Float_32_Div_altfp_div_csa_ovb
	  PORT MAP ( 
		dataa => srt_adjust_w,
		datab => value_one_w,
		result => wire_altfp_div_csa27_result
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_next_special_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN divider_next_special_dffe <= divider_next_w13c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN Rk_remainder_special_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN Rk_remainder_special_dffe <= Rk_next_w13c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe0c <= ( rom_reg_dffe0c(47 DOWNTO 0) & rom_out_w0c(1 DOWNTO 0));
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe10c <= ( rom_reg_dffe10c(11 DOWNTO 0) & rom_out_w10c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe11c <= ( rom_reg_dffe11c(5 DOWNTO 0) & rom_out_w11c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe12c <= ( rom_out_w12c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe1c <= ( rom_reg_dffe1c(65 DOWNTO 0) & rom_out_w1c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe2c <= ( rom_reg_dffe2c(59 DOWNTO 0) & rom_out_w2c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe3c <= ( rom_reg_dffe3c(53 DOWNTO 0) & rom_out_w3c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe4c <= ( rom_reg_dffe4c(47 DOWNTO 0) & rom_out_w4c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe5c <= ( rom_reg_dffe5c(41 DOWNTO 0) & rom_out_w5c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe6c <= ( rom_reg_dffe6c(35 DOWNTO 0) & rom_out_w6c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe7c <= ( rom_reg_dffe7c(29 DOWNTO 0) & rom_out_w7c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe8c <= ( rom_reg_dffe8c(23 DOWNTO 0) & rom_out_w8c);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rom_reg_dffe9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clken = '1') THEN rom_reg_dffe9c <= ( rom_reg_dffe9c(17 DOWNTO 0) & rom_out_w9c);
			END IF;
		END IF;
	END PROCESS;
	srt_block_int11 :  Float_32_Div_srt_block_int_sfk
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_w,
		divider_reg => wire_srt_block_int11_divider_reg,
		Rk => Rk_w,
		Rk_next => wire_srt_block_int11_Rk_next,
		rom => wire_srt_block_int11_rom
	  );
	srt_block_int12 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w0c,
		divider_reg => wire_srt_block_int12_divider_reg,
		Rk => Rk_next_w0c,
		Rk_next => wire_srt_block_int12_Rk_next,
		rom => wire_srt_block_int12_rom
	  );
	srt_block_int13 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w1c,
		divider_reg => wire_srt_block_int13_divider_reg,
		Rk => Rk_next_w1c,
		Rk_next => wire_srt_block_int13_Rk_next,
		rom => wire_srt_block_int13_rom
	  );
	srt_block_int14 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w2c,
		divider_reg => wire_srt_block_int14_divider_reg,
		Rk => Rk_next_w2c,
		Rk_next => wire_srt_block_int14_Rk_next,
		rom => wire_srt_block_int14_rom
	  );
	srt_block_int15 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w3c,
		divider_reg => wire_srt_block_int15_divider_reg,
		Rk => Rk_next_w3c,
		Rk_next => wire_srt_block_int15_Rk_next,
		rom => wire_srt_block_int15_rom
	  );
	srt_block_int16 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w4c,
		divider_reg => wire_srt_block_int16_divider_reg,
		Rk => Rk_next_w4c,
		Rk_next => wire_srt_block_int16_Rk_next,
		rom => wire_srt_block_int16_rom
	  );
	srt_block_int17 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w5c,
		divider_reg => wire_srt_block_int17_divider_reg,
		Rk => Rk_next_w5c,
		Rk_next => wire_srt_block_int17_Rk_next,
		rom => wire_srt_block_int17_rom
	  );
	srt_block_int18 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w6c,
		divider_reg => wire_srt_block_int18_divider_reg,
		Rk => Rk_next_w6c,
		Rk_next => wire_srt_block_int18_Rk_next,
		rom => wire_srt_block_int18_rom
	  );
	srt_block_int19 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w7c,
		divider_reg => wire_srt_block_int19_divider_reg,
		Rk => Rk_next_w7c,
		Rk_next => wire_srt_block_int19_Rk_next,
		rom => wire_srt_block_int19_rom
	  );
	srt_block_int20 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w8c,
		divider_reg => wire_srt_block_int20_divider_reg,
		Rk => Rk_next_w8c,
		Rk_next => wire_srt_block_int20_Rk_next,
		rom => wire_srt_block_int20_rom
	  );
	srt_block_int21 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w9c,
		divider_reg => wire_srt_block_int21_divider_reg,
		Rk => Rk_next_w9c,
		Rk_next => wire_srt_block_int21_Rk_next,
		rom => wire_srt_block_int21_rom
	  );
	srt_block_int22 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w10c,
		divider_reg => wire_srt_block_int22_divider_reg,
		Rk => Rk_next_w10c,
		Rk_next => wire_srt_block_int22_Rk_next,
		rom => wire_srt_block_int22_rom
	  );
	srt_block_int23 :  Float_32_Div_srt_block_int_4ik
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w11c,
		divider_reg => wire_srt_block_int23_divider_reg,
		Rk => Rk_next_w11c,
		Rk_next => wire_srt_block_int23_Rk_next,
		rom => wire_srt_block_int23_rom
	  );
	srt_block_int24 :  Float_32_Div_srt_block_int_bck
	  PORT MAP ( 
		aclr => aclr,
		clken => clken,
		clock => clock,
		divider => divider_next_w12c,
		divider_reg => wire_srt_block_int24_divider_reg,
		Rk => Rk_next_w12c,
		Rk_next => wire_srt_block_int24_Rk_next,
		rom => wire_srt_block_int24_rom
	  );

 END RTL; --Float_32_Div_altfp_div_srt_ext_14f

 LIBRARY lpm;
 USE lpm.all;

--synthesis_resources = lpm_add_sub 21 lpm_compare 62 lpm_mux 28 reg 2690 
 LIBRARY ieee;
 USE ieee.std_logic_1164.all;

 ENTITY  Float_32_Div_altfp_div_01j IS 
	 PORT 
	 ( 
		 clock	:	IN  STD_LOGIC;
		 dataa	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 datab	:	IN  STD_LOGIC_VECTOR (31 DOWNTO 0);
		 division_by_zero	:	OUT  STD_LOGIC;
		 result	:	OUT  STD_LOGIC_VECTOR (31 DOWNTO 0)
	 ); 
 END Float_32_Div_altfp_div_01j;

 ARCHITECTURE RTL OF Float_32_Div_altfp_div_01j IS

	 SIGNAL  wire_altfp_div_csa8_cout	:	STD_LOGIC;
	 SIGNAL  wire_altfp_div_csa8_result	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_divider	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_quotient	:	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  wire_altfp_div_srt_ext1_remain	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL	 and_or_dffe	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_dffe1a	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_dffe3a	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline0c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline10c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline11c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline12c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline13c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline14c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline15c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline16c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline17c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline18c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline19c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline1c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline20c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline21c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline22c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline23c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline24c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline25c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline26c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline27c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline2c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline3c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline4c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline5c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline6c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline7c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline8c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 and_or_pipeline9c	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 bias_addition_overf_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_bias_addition_overf_dffe_w_lg_q781w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 divider_pipe1a	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 division_by_zero_port_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_a_and_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_a_b_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_a_dffe	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_a_or_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_a_or_dffe_w_lg_q629w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exp_b_and_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_b_dffe	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_b_or_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_exp_b_or_dffe_w_lg_q632w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 exp_dffe1a	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_dffe2a	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline0c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline10c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline11c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline12c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline13c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline14c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline15c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline16c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline17c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline18c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline19c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline1c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline20c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline21c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline22c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline23c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline24c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline25c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline26c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline2c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline3c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline4c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline5c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline6c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline7c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline8c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_pipeline9c	:	STD_LOGIC_VECTOR(8 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 exp_res_pipe3	:	STD_LOGIC_VECTOR(7 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 implied_bit	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 implied_bit2a	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_a_and_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_a_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_a_or_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_a_or_dffe_w_lg_q635w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_b_and_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_b_dffe	:	STD_LOGIC_VECTOR(22 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 man_b_or_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_man_b_or_dffe_w_lg_q638w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL	 man_res_pipe3	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 quotient_pipe1a	:	STD_LOGIC_VECTOR(27 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 remainder_pipe1a	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 result_output_dffe	:	STD_LOGIC_VECTOR(31 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rnd_overflow_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 rnded_man_pipe2a	:	STD_LOGIC_VECTOR(23 DOWNTO 0)
	 -- synopsys translate_off
	  := (OTHERS => '0')
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_a_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_b_dffe	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline0c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline10c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline11c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline12c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline13c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline14c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline15c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline16c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline17c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline18c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline19c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline1c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline20c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline21c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline22c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline23c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline24c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline25c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline26c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline27c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline2c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline3c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline4c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline5c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline6c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline7c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline8c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_div_pipeline9c	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe1a	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe2a	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL	 sign_pipe3a	:	STD_LOGIC
	 -- synopsys translate_off
	  := '0'
	 -- synopsys translate_on
	 ;
	 SIGNAL  wire_add_sub10_overflow	:	STD_LOGIC;
	 SIGNAL  wire_add_sub10_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_add_sub9_result	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_cmpr2_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr2_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr3_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr4_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr5_ageb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr6_aeb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr6_agb	:	STD_LOGIC;
	 SIGNAL  wire_cmpr7_ageb	:	STD_LOGIC;
	 SIGNAL  wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w524w525w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w522w523w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_guard_bit_dffe1a_w446w447w448w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w481w482w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w479w480w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bias_addition_overf_w519w520w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux1_exp_s1a476w477w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux1_exp_s1a473w474w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bias_addition_overf_w521w524w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_bias_addition_overf_w521w522w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0329w333w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0329w330w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0329w337w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0329w335w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0329w353w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0339w343w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0339w340w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0339w347w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0339w345w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0339w361w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_a_b_w487w488w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_guard_bit_dffe1a_w446w447w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_infinite_w800w801w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux1_exp_s1a478w481w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux1_exp_s1a478w479w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_mux_zero_non_zero_S0590w591w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_nan_w780w808w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w621w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w624w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_quo_msb_m1_w380w436w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_quo_msb_m1_w380w381w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_quo_msb_m1_w380w439w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_quo_msb_m1_w380w442w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_rnd_overflow457w458w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_zero_w804w805w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_bias_addition_overf_w519w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dataa_S0354w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_datab_S0362w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_b_w486w	:	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_non_zero_w643w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_b_non_zero_w652w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_infi_bus_w586w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinite_w802w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux1_exp_s1a476w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux1_exp_s1a473w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_zero_non_zero_S0592w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_w809w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_exp_res_int2_or_res_w625w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_exp_res_int2_or_res_w622w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_lg_quo_msb_m1_w382w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w_lg_rnd_overflow459w	:	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  wire_w411w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_w806w	:	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range26w28w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range29w30w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range31w32w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range33w34w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range35w36w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range37w38w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_and_w_range39w40w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range67w69w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range70w71w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range72w73w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range74w75w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range76w77w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range78w79w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_and_w_range80w81w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range492w495w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range496w498w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range499w501w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range502w504w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range505w507w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range508w510w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_bias_and_w_range511w513w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range680w683w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range684w686w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range687w689w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range690w692w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range693w695w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range696w698w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_and_w_range699w701w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range153w155w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range174w175w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range176w177w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range178w179w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range180w181w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range182w183w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range184w185w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range186w187w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range188w189w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range190w191w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range192w193w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range156w157w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range194w195w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range196w197w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range158w159w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range160w161w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range162w163w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range164w165w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range166w167w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range168w169w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range170w171w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_and_w_range172w173w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range269w271w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range290w291w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range292w293w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range294w295w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range296w297w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range298w299w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range300w301w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range302w303w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range304w305w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range306w307w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range308w309w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range272w273w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range310w311w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range312w313w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range274w275w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range276w277w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range278w279w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range280w281w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range282w283w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range284w285w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range286w287w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_and_w_range288w289w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range562w565w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range566w568w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range569w571w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range572w574w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range575w577w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range578w580w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_infi_and_w_range581w583w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_bias_addition_overf_w521w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_dataa_S0329w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_datab_S0339w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_b_w487w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_one_w640w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_a_or_msb_w325w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_b_one_w649w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_b_or_msb_w327w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_sign_w516w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_guard_bit_dffe1a_w446w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infi_combi_w779w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_infinite_w800w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux1_exp_s0a475w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux1_exp_s1a478w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_mux_zero_non_zero_S0590w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_nan_w780w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_not_exp_res_int2_or_res_w620w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_quo_msb_m1_w380w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_rnd_overflow457w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_dataa_w775w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_zero_w804w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range772w773w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_dataa_S0354w355w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_datab_S0362w363w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_exp_zero_bus_w587w588w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_a_zero_w641w642w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_lg_man_b_zero_w650w651w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_exp_zero_bus_w587w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_a_zero_w641w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_man_b_zero_w650w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w412w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range3w6w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range7w9w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range10w12w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range13w15w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range16w18w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range19w21w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_a_or_w_range22w24w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range44w47w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range48w50w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range51w53w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range54w56w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range57w59w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range60w62w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_b_or_w_range63w65w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_higher_or_range531w534w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range596w599w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range600w602w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range603w605w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range606w608w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range609w611w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range612w614w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_exp_res_int2_or_w_range615w617w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range85w88w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range116w118w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range119w121w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range122w124w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range125w127w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range128w130w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range131w133w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range134w136w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range137w139w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range140w142w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range143w145w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range89w91w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range146w148w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range149w151w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range92w94w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range95w97w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range98w100w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range101w103w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range104w106w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range107w109w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range110w112w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_a_or_w_range113w115w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range201w204w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range232w234w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range235w237w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range238w240w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range241w243w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range244w246w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range247w249w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range250w252w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range253w255w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range256w258w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range259w261w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range205w207w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range262w264w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range265w267w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range208w210w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range211w213w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range214w216w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range217w219w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range220w222w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range223w225w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range226w228w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_b_or_w_range229w231w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range705w708w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range736w738w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range739w741w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range742w744w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range745w747w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range748w750w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range751w753w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range754w756w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range757w759w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range760w762w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range763w765w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range709w711w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range766w768w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range769w771w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range712w714w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range715w717w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range718w720w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range721w723w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range724w726w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range727w729w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range730w732w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_man_res_or_w_range733w735w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range537w540w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range541w543w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range544w546w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range547w549w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range550w552w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range553w555w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_norm_zero_or_w_range556w558w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_lg_w_sticky_bit_quo_msb_m1_or_range388w391w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  aclr	:	STD_LOGIC;
	 SIGNAL  add_1_dataa_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  add_1_datab_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  add_1_w :	STD_LOGIC;
	 SIGNAL  add_one_process_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  and_or_dffe1a_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  and_or_dffe3a_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  and_or_dffe_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  and_or_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  and_or_pipeline_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bias_add_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  bias_addition_overf_w :	STD_LOGIC;
	 SIGNAL  bias_addition_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  bias_value_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  checked_quotient_dffe1a_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  checked_quotient_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  clk_en	:	STD_LOGIC;
	 SIGNAL  dataa_exp_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  dataa_int :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  dataa_man_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  dataa_S0 :	STD_LOGIC;
	 SIGNAL  datab_exp_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  datab_int :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  datab_man_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  datab_S0 :	STD_LOGIC;
	 SIGNAL  divider_srt_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  division_by_w :	STD_LOGIC;
	 SIGNAL  exp_a_and_msb2_w :	STD_LOGIC;
	 SIGNAL  exp_a_and_msb_w :	STD_LOGIC;
	 SIGNAL  exp_a_and_mux_w :	STD_LOGIC;
	 SIGNAL  exp_a_and_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_b_w :	STD_LOGIC;
	 SIGNAL  exp_a_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_non_zero_w :	STD_LOGIC;
	 SIGNAL  exp_a_one_w :	STD_LOGIC;
	 SIGNAL  exp_a_or_msb2_w :	STD_LOGIC;
	 SIGNAL  exp_a_or_msb_w :	STD_LOGIC;
	 SIGNAL  exp_a_or_mux_w :	STD_LOGIC;
	 SIGNAL  exp_a_or_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_a_zero_w :	STD_LOGIC;
	 SIGNAL  exp_b_and_msb2_w :	STD_LOGIC;
	 SIGNAL  exp_b_and_msb_w :	STD_LOGIC;
	 SIGNAL  exp_b_and_mux_w :	STD_LOGIC;
	 SIGNAL  exp_b_and_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_non_zero_w :	STD_LOGIC;
	 SIGNAL  exp_b_one_w :	STD_LOGIC;
	 SIGNAL  exp_b_or_msb2_w :	STD_LOGIC;
	 SIGNAL  exp_b_or_msb_w :	STD_LOGIC;
	 SIGNAL  exp_b_or_mux_w :	STD_LOGIC;
	 SIGNAL  exp_b_or_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_b_zero_w :	STD_LOGIC;
	 SIGNAL  exp_bias_and_res_w :	STD_LOGIC;
	 SIGNAL  exp_bias_and_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_bias_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_dffe1a_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_dffe2a_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_exc_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_exc_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_higher_bit :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_higher_or :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  exp_infi_bus_w :	STD_LOGIC;
	 SIGNAL  exp_man_and_or_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_or_result_w :	STD_LOGIC;
	 SIGNAL  exp_pipeline_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_res_and_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_int2_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_int2_or_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_int2_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_int_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_res_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  exp_sign_w :	STD_LOGIC;
	 SIGNAL  exp_sub_a_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_b_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_sub_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  exp_zero_bus_w :	STD_LOGIC;
	 SIGNAL  guard_bit_dffe1a_w :	STD_LOGIC;
	 SIGNAL  guard_bit_quo_msb_m1 :	STD_LOGIC;
	 SIGNAL  guard_bit_quo_msb_m2 :	STD_LOGIC;
	 SIGNAL  guard_bit_w :	STD_LOGIC;
	 SIGNAL  infi_combi_w :	STD_LOGIC;
	 SIGNAL  infi_dataa_w :	STD_LOGIC;
	 SIGNAL  infi_datab_w :	STD_LOGIC;
	 SIGNAL  infi_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  infinite_int_w :	STD_LOGIC;
	 SIGNAL  infinite_w :	STD_LOGIC;
	 SIGNAL  man_24_zeros_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_a_and_msb2_w :	STD_LOGIC;
	 SIGNAL  man_a_and_msb_w :	STD_LOGIC;
	 SIGNAL  man_a_and_mux_w :	STD_LOGIC;
	 SIGNAL  man_a_and_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_int_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_non_zero_w :	STD_LOGIC;
	 SIGNAL  man_a_one_w :	STD_LOGIC;
	 SIGNAL  man_a_or_msb2_w :	STD_LOGIC;
	 SIGNAL  man_a_or_msb_w :	STD_LOGIC;
	 SIGNAL  man_a_or_mux_w :	STD_LOGIC;
	 SIGNAL  man_a_or_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_a_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_a_zero_w :	STD_LOGIC;
	 SIGNAL  man_b_and_msb2_w :	STD_LOGIC;
	 SIGNAL  man_b_and_msb_w :	STD_LOGIC;
	 SIGNAL  man_b_and_mux_w :	STD_LOGIC;
	 SIGNAL  man_b_and_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_int_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_non_zero_w :	STD_LOGIC;
	 SIGNAL  man_b_one_w :	STD_LOGIC;
	 SIGNAL  man_b_or_msb2_w :	STD_LOGIC;
	 SIGNAL  man_b_or_msb_w :	STD_LOGIC;
	 SIGNAL  man_b_or_mux_w :	STD_LOGIC;
	 SIGNAL  man_b_or_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_b_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_b_zero_w :	STD_LOGIC;
	 SIGNAL  man_exc_nan_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_exc_zeros_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_bus_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_int2_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_res_int_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  man_res_or_w :	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  man_res_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  mux1_exp_s0a :	STD_LOGIC;
	 SIGNAL  mux1_exp_s1a :	STD_LOGIC;
	 SIGNAL  mux_1_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mux_2_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mux_3_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  mux_zero_non_zero_S0 :	STD_LOGIC;
	 SIGNAL  mux_zero_non_zero_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  nan_dataa_w :	STD_LOGIC;
	 SIGNAL  nan_datab_w :	STD_LOGIC;
	 SIGNAL  nan_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  nan_w :	STD_LOGIC;
	 SIGNAL  norm_dataa_w :	STD_LOGIC;
	 SIGNAL  norm_datab_w :	STD_LOGIC;
	 SIGNAL  norm_infi_and_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  norm_infi_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  norm_res_int_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  norm_zero_bus_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  norm_zero_or_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  not_bias_addition_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  not_exp_res_int2_or_res_w :	STD_LOGIC;
	 SIGNAL  overflow_int_w :	STD_LOGIC;
	 SIGNAL  overflow_man_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  overflow_ones_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  quo_msb_m1_compare_dataa :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  quo_msb_m1_compare_datab :	STD_LOGIC_VECTOR (52 DOWNTO 0);
	 SIGNAL  quo_msb_m1_compare_w :	STD_LOGIC;
	 SIGNAL  quo_msb_m1_w :	STD_LOGIC;
	 SIGNAL  quo_msb_m2_compare_dataa :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  quo_msb_m2_compare_datab :	STD_LOGIC_VECTOR (53 DOWNTO 0);
	 SIGNAL  quo_msb_m2_compare_w :	STD_LOGIC;
	 SIGNAL  quotient_msb_m1_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  quotient_msb_m2_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  quotient_w :	STD_LOGIC_VECTOR (27 DOWNTO 0);
	 SIGNAL  remainder_srt_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  res_rnded_man_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  rnd_add_overf_w :	STD_LOGIC;
	 SIGNAL  rnd_overflow :	STD_LOGIC;
	 SIGNAL  rnded_man_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  round_bit_dffe1a_w :	STD_LOGIC;
	 SIGNAL  round_bit_quo_msb_m1 :	STD_LOGIC;
	 SIGNAL  round_bit_quo_msb_m2 :	STD_LOGIC;
	 SIGNAL  round_bit_w :	STD_LOGIC;
	 SIGNAL  sign_a_w :	STD_LOGIC;
	 SIGNAL  sign_b_w :	STD_LOGIC;
	 SIGNAL  sign_div :	STD_LOGIC;
	 SIGNAL  sign_div_pipeline_w :	STD_LOGIC;
	 SIGNAL  sign_exc_bit_w :	STD_LOGIC;
	 SIGNAL  signed_N_exp_h_or :	STD_LOGIC;
	 SIGNAL  sticky_bit_dffe1a_w :	STD_LOGIC;
	 SIGNAL  sticky_bit_quo_msb_m1 :	STD_LOGIC;
	 SIGNAL  sticky_bit_quo_msb_m1_bit :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  sticky_bit_quo_msb_m1_or :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  sticky_bit_quo_msb_m1_tmp :	STD_LOGIC_VECTOR (1 DOWNTO 0);
	 SIGNAL  sticky_bit_quo_msb_m2 :	STD_LOGIC;
	 SIGNAL  sticky_bit_quo_msb_m2_bit :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sticky_bit_quo_msb_m2_or :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sticky_bit_quo_msb_m2_tmp :	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  sticky_bit_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_lower_lower_ageb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_lower_upper_aeb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_lower_upper_agb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_upper_lower_aeb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_upper_lower_agb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_upper_upper_aeb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m1_comparator_upper_upper_agb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m2_comparator_lower_ageb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m2_comparator_upper_aeb_w :	STD_LOGIC;
	 SIGNAL  sticky_quo_msb_m2_comparator_upper_agb_w :	STD_LOGIC;
	 SIGNAL  underflow_zeros_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  value_add_1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_minus_1_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_normal_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  value_zero_w :	STD_LOGIC_VECTOR (8 DOWNTO 0);
	 SIGNAL  zero_bit_23_w :	STD_LOGIC_VECTOR (23 DOWNTO 0);
	 SIGNAL  zero_bit_31_w :	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  zero_bit_8_w :	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  zero_bit_w :	STD_LOGIC;
	 SIGNAL  zero_dataa_w :	STD_LOGIC;
	 SIGNAL  zero_datab_w :	STD_LOGIC;
	 SIGNAL  zero_res_w :	STD_LOGIC_VECTOR (31 DOWNTO 0);
	 SIGNAL  zero_w :	STD_LOGIC;
	 SIGNAL  wire_w_dataa_range352w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_dataa_int_range366w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_dataa_int_range365w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_datab_range360w	:	STD_LOGIC_VECTOR (30 DOWNTO 0);
	 SIGNAL  wire_w_datab_int_range368w	:	STD_LOGIC_VECTOR (22 DOWNTO 0);
	 SIGNAL  wire_w_datab_int_range367w	:	STD_LOGIC_VECTOR (7 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range26w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range29w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range31w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range33w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range35w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range37w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_and_w_range39w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range5w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range8w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range11w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range14w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range17w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range20w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_bus_w_range23w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range3w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range7w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range10w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range13w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range16w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range19w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_a_or_w_range22w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range67w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range70w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range72w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range74w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range76w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range78w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_and_w_range80w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range46w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range49w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range52w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range55w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range58w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range61w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_bus_w_range64w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range44w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range48w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range51w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range54w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range57w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range60w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_b_or_w_range63w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range492w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range496w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range499w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range502w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range505w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range508w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_and_w_range511w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range494w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range497w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range500w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range503w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range506w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range509w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_bias_bus_w_range512w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_higher_bit_range533w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_higher_or_range531w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range680w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range684w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range687w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range690w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range693w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range696w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range699w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_and_w_range702w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range682w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range685w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range688w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range691w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range694w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range697w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_bus_w_range700w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range598w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range601w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range604w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range607w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range610w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range613w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_bus_w_range616w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range596w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range600w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range603w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range606w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range609w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range612w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_exp_res_int2_or_w_range615w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range153w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range174w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range176w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range178w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range180w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range182w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range184w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range186w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range188w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range190w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range192w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range156w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range194w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range196w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range158w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range160w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range162w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range164w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range166w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range168w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range170w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_and_w_range172w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range114w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range117w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range120w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range123w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range126w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range129w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range132w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range135w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range138w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range141w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range87w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range144w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range147w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range150w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range90w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range93w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range96w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range99w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range102w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range105w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range108w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_bus_w_range111w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range85w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range116w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range119w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range122w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range125w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range128w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range131w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range134w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range137w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range140w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range143w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range89w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range146w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range149w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range92w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range95w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range98w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range101w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range104w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range107w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range110w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_a_or_w_range113w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range269w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range290w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range292w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range294w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range296w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range298w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range300w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range302w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range304w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range306w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range308w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range272w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range310w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range312w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range274w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range276w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range278w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range280w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range282w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range284w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range286w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_and_w_range288w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range230w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range233w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range236w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range239w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range242w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range245w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range248w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range251w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range254w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range257w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range203w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range260w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range263w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range266w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range206w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range209w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range212w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range215w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range218w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range221w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range224w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_bus_w_range227w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range201w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range232w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range235w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range238w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range241w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range244w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range247w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range250w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range253w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range256w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range259w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range205w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range262w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range265w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range208w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range211w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range214w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range217w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range220w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range223w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range226w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_b_or_w_range229w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range734w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range737w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range740w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range743w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range746w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range749w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range752w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range755w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range758w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range761w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range707w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range764w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range767w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range770w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range710w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range713w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range716w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range719w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range722w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range725w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range728w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_bus_w_range731w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range705w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range736w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range739w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range742w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range745w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range748w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range751w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range754w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range757w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range760w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range763w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range709w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range766w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range769w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range772w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range712w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range715w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range718w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range721w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range724w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range727w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range730w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_man_res_or_w_range733w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range562w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range566w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range569w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range572w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range575w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range578w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_and_w_range581w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range564w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range567w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range570w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range573w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range576w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range579w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_infi_bus_w_range582w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range539w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range542w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range545w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range548w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range551w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range554w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_bus_w_range557w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range537w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range541w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range544w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range547w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range550w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range553w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_norm_zero_or_w_range556w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_quo_msb_m1_bit_range390w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 SIGNAL  wire_w_sticky_bit_quo_msb_m1_or_range388w	:	STD_LOGIC_VECTOR (0 DOWNTO 0);
	 COMPONENT  Float_32_Div_altfp_div_csa_gvc
	 PORT
	 ( 
		cin	:	IN  STD_LOGIC := '0';
		cout	:	OUT  STD_LOGIC;
		dataa	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0) := (OTHERS => '0');
		result	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  Float_32_Div_altfp_div_srt_ext_14f
	 PORT
	 ( 
		aclr	:	IN  STD_LOGIC := '0';
		clken	:	IN  STD_LOGIC := '1';
		clock	:	IN  STD_LOGIC := '0';
		denom	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		divider	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0);
		numer	:	IN  STD_LOGIC_VECTOR(23 DOWNTO 0);
		quotient	:	OUT  STD_LOGIC_VECTOR(27 DOWNTO 0);
		remain	:	OUT  STD_LOGIC_VECTOR(23 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_add_sub
	 GENERIC 
	 (
		LPM_DIRECTION	:	STRING := "DEFAULT";
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "SIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_add_sub"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		add_sub	:	IN STD_LOGIC := '1';
		cin	:	IN STD_LOGIC := 'Z';
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		cout	:	OUT STD_LOGIC;
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		overflow	:	OUT STD_LOGIC;
		result	:	OUT STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0)
	 ); 
	 END COMPONENT;
	 COMPONENT  lpm_compare
	 GENERIC 
	 (
		LPM_PIPELINE	:	NATURAL := 0;
		LPM_REPRESENTATION	:	STRING := "UNSIGNED";
		LPM_WIDTH	:	NATURAL;
		lpm_hint	:	STRING := "UNUSED";
		lpm_type	:	STRING := "lpm_compare"
	 );
	 PORT
	 ( 
		aclr	:	IN STD_LOGIC := '0';
		aeb	:	OUT STD_LOGIC;
		agb	:	OUT STD_LOGIC;
		ageb	:	OUT STD_LOGIC;
		alb	:	OUT STD_LOGIC;
		aleb	:	OUT STD_LOGIC;
		aneb	:	OUT STD_LOGIC;
		clken	:	IN STD_LOGIC := '1';
		clock	:	IN STD_LOGIC := '0';
		dataa	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0');
		datab	:	IN STD_LOGIC_VECTOR(LPM_WIDTH-1 DOWNTO 0) := (OTHERS => '0')
	 ); 
	 END COMPONENT;
 BEGIN

	loop73 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w524w525w(i) <= wire_w_lg_w_lg_bias_addition_overf_w521w524w(0) AND bias_addition_w(i);
	END GENERATE loop73;
	loop74 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w522w523w(i) <= wire_w_lg_w_lg_bias_addition_overf_w521w522w(0) AND underflow_zeros_w(i);
	END GENERATE loop74;
	wire_w_lg_w_lg_w_lg_guard_bit_dffe1a_w446w447w448w(0) <= wire_w_lg_w_lg_guard_bit_dffe1a_w446w447w(0) AND sticky_bit_dffe1a_w;
	loop75 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w481w482w(i) <= wire_w_lg_w_lg_mux1_exp_s1a478w481w(0) AND value_minus_1_w(i);
	END GENERATE loop75;
	loop76 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w479w480w(i) <= wire_w_lg_w_lg_mux1_exp_s1a478w479w(0) AND value_normal_w(i);
	END GENERATE loop76;
	loop77 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_bias_addition_overf_w519w520w(i) <= wire_w_lg_bias_addition_overf_w519w(0) AND overflow_ones_w(i);
	END GENERATE loop77;
	loop78 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_mux1_exp_s1a476w477w(i) <= wire_w_lg_mux1_exp_s1a476w(0) AND value_normal_w(i);
	END GENERATE loop78;
	loop79 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_mux1_exp_s1a473w474w(i) <= wire_w_lg_mux1_exp_s1a473w(0) AND value_add_1_w(i);
	END GENERATE loop79;
	wire_w_lg_w_lg_bias_addition_overf_w521w524w(0) <= wire_w_lg_bias_addition_overf_w521w(0) AND wire_w_lg_exp_sign_w516w(0);
	wire_w_lg_w_lg_bias_addition_overf_w521w522w(0) <= wire_w_lg_bias_addition_overf_w521w(0) AND exp_sign_w;
	wire_w_lg_w_lg_dataa_S0329w333w(0) <= wire_w_lg_dataa_S0329w(0) AND exp_a_and_msb_w;
	wire_w_lg_w_lg_dataa_S0329w330w(0) <= wire_w_lg_dataa_S0329w(0) AND exp_a_or_msb_w;
	wire_w_lg_w_lg_dataa_S0329w337w(0) <= wire_w_lg_dataa_S0329w(0) AND man_a_and_msb_w;
	wire_w_lg_w_lg_dataa_S0329w335w(0) <= wire_w_lg_dataa_S0329w(0) AND man_a_or_msb_w;
	loop80 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_dataa_S0329w353w(i) <= wire_w_lg_dataa_S0329w(0) AND wire_w_dataa_range352w(i);
	END GENERATE loop80;
	wire_w_lg_w_lg_datab_S0339w343w(0) <= wire_w_lg_datab_S0339w(0) AND exp_b_and_msb_w;
	wire_w_lg_w_lg_datab_S0339w340w(0) <= wire_w_lg_datab_S0339w(0) AND exp_b_or_msb_w;
	wire_w_lg_w_lg_datab_S0339w347w(0) <= wire_w_lg_datab_S0339w(0) AND man_b_and_msb_w;
	wire_w_lg_w_lg_datab_S0339w345w(0) <= wire_w_lg_datab_S0339w(0) AND man_b_or_msb_w;
	loop81 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_datab_S0339w361w(i) <= wire_w_lg_datab_S0339w(0) AND wire_w_datab_range360w(i);
	END GENERATE loop81;
	loop82 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_w_lg_exp_a_b_w487w488w(i) <= wire_w_lg_exp_a_b_w487w(0) AND value_zero_w(i);
	END GENERATE loop82;
	wire_w_lg_w_lg_guard_bit_dffe1a_w446w447w(0) <= wire_w_lg_guard_bit_dffe1a_w446w(0) AND round_bit_dffe1a_w;
	loop83 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_infinite_w800w801w(i) <= wire_w_lg_infinite_w800w(0) AND norm_res_int_w(i);
	END GENERATE loop83;
	wire_w_lg_w_lg_mux1_exp_s1a478w481w(0) <= wire_w_lg_mux1_exp_s1a478w(0) AND wire_w_lg_mux1_exp_s0a475w(0);
	wire_w_lg_w_lg_mux1_exp_s1a478w479w(0) <= wire_w_lg_mux1_exp_s1a478w(0) AND mux1_exp_s0a;
	loop84 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_w_lg_mux_zero_non_zero_S0590w591w(i) <= wire_w_lg_mux_zero_non_zero_S0590w(0) AND res_rnded_man_w(i);
	END GENERATE loop84;
	loop85 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_nan_w780w808w(i) <= wire_w_lg_nan_w780w(0) AND mux_2_res_w(i);
	END GENERATE loop85;
	loop86 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w621w(i) <= wire_w_lg_not_exp_res_int2_or_res_w620w(0) AND exp_res_int2_w(i);
	END GENERATE loop86;
	loop87 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w624w(i) <= wire_w_lg_not_exp_res_int2_or_res_w620w(0) AND man_res_int2_w(i);
	END GENERATE loop87;
	wire_w_lg_w_lg_quo_msb_m1_w380w436w(0) <= wire_w_lg_quo_msb_m1_w380w(0) AND guard_bit_quo_msb_m2;
	loop88 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_w_lg_quo_msb_m1_w380w381w(i) <= wire_w_lg_quo_msb_m1_w380w(0) AND quotient_msb_m2_w(i);
	END GENERATE loop88;
	wire_w_lg_w_lg_quo_msb_m1_w380w439w(0) <= wire_w_lg_quo_msb_m1_w380w(0) AND round_bit_quo_msb_m2;
	wire_w_lg_w_lg_quo_msb_m1_w380w442w(0) <= wire_w_lg_quo_msb_m1_w380w(0) AND sticky_bit_quo_msb_m2;
	loop89 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_w_lg_rnd_overflow457w458w(i) <= wire_w_lg_rnd_overflow457w(0) AND add_one_process_w(i);
	END GENERATE loop89;
	loop90 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_w_lg_zero_w804w805w(i) <= wire_w_lg_zero_w804w(0) AND mux_1_res_w(i);
	END GENERATE loop90;
	wire_w_lg_bias_addition_overf_w519w(0) <= bias_addition_overf_w AND wire_w_lg_exp_sign_w516w(0);
	loop91 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_dataa_S0354w(i) <= dataa_S0 AND zero_bit_31_w(i);
	END GENERATE loop91;
	loop92 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_datab_S0362w(i) <= datab_S0 AND zero_bit_31_w(i);
	END GENERATE loop92;
	loop93 : FOR i IN 0 TO 8 GENERATE 
		wire_w_lg_exp_a_b_w486w(i) <= exp_a_b_w AND bias_value_w(i);
	END GENERATE loop93;
	wire_w_lg_exp_a_non_zero_w643w(0) <= exp_a_non_zero_w AND wire_w_lg_w_lg_man_a_zero_w641w642w(0);
	wire_w_lg_exp_b_non_zero_w652w(0) <= exp_b_non_zero_w AND wire_w_lg_w_lg_man_b_zero_w650w651w(0);
	wire_w_lg_exp_infi_bus_w586w(0) <= exp_infi_bus_w AND wire_w_lg_exp_sign_w516w(0);
	loop94 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_infinite_w802w(i) <= infinite_w AND infi_res_w(i);
	END GENERATE loop94;
	wire_w_lg_mux1_exp_s1a476w(0) <= mux1_exp_s1a AND wire_w_lg_mux1_exp_s0a475w(0);
	wire_w_lg_mux1_exp_s1a473w(0) <= mux1_exp_s1a AND mux1_exp_s0a;
	loop95 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_mux_zero_non_zero_S0592w(i) <= mux_zero_non_zero_S0 AND man_24_zeros_w(i);
	END GENERATE loop95;
	loop96 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_nan_w809w(i) <= nan_w AND nan_res_w(i);
	END GENERATE loop96;
	loop97 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_not_exp_res_int2_or_res_w625w(i) <= not_exp_res_int2_or_res_w AND zero_bit_23_w(i);
	END GENERATE loop97;
	loop98 : FOR i IN 0 TO 7 GENERATE 
		wire_w_lg_not_exp_res_int2_or_res_w622w(i) <= not_exp_res_int2_or_res_w AND zero_bit_8_w(i);
	END GENERATE loop98;
	loop99 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_quo_msb_m1_w382w(i) <= quo_msb_m1_w AND quotient_msb_m1_w(i);
	END GENERATE loop99;
	loop100 : FOR i IN 0 TO 23 GENERATE 
		wire_w_lg_rnd_overflow459w(i) <= rnd_overflow AND overflow_man_w(i);
	END GENERATE loop100;
	wire_w411w(0) <= sticky_quo_msb_m1_comparator_upper_upper_aeb_w AND sticky_quo_msb_m1_comparator_upper_lower_agb_w;
	loop101 : FOR i IN 0 TO 31 GENERATE 
		wire_w_lg_zero_w806w(i) <= zero_w AND zero_res_w(i);
	END GENERATE loop101;
	wire_w_lg_w_exp_a_and_w_range26w28w(0) <= wire_w_exp_a_and_w_range26w(0) AND wire_w_exp_a_bus_w_range5w(0);
	wire_w_lg_w_exp_a_and_w_range29w30w(0) <= wire_w_exp_a_and_w_range29w(0) AND wire_w_exp_a_bus_w_range8w(0);
	wire_w_lg_w_exp_a_and_w_range31w32w(0) <= wire_w_exp_a_and_w_range31w(0) AND wire_w_exp_a_bus_w_range11w(0);
	wire_w_lg_w_exp_a_and_w_range33w34w(0) <= wire_w_exp_a_and_w_range33w(0) AND wire_w_exp_a_bus_w_range14w(0);
	wire_w_lg_w_exp_a_and_w_range35w36w(0) <= wire_w_exp_a_and_w_range35w(0) AND wire_w_exp_a_bus_w_range17w(0);
	wire_w_lg_w_exp_a_and_w_range37w38w(0) <= wire_w_exp_a_and_w_range37w(0) AND wire_w_exp_a_bus_w_range20w(0);
	wire_w_lg_w_exp_a_and_w_range39w40w(0) <= wire_w_exp_a_and_w_range39w(0) AND wire_w_exp_a_bus_w_range23w(0);
	wire_w_lg_w_exp_b_and_w_range67w69w(0) <= wire_w_exp_b_and_w_range67w(0) AND wire_w_exp_b_bus_w_range46w(0);
	wire_w_lg_w_exp_b_and_w_range70w71w(0) <= wire_w_exp_b_and_w_range70w(0) AND wire_w_exp_b_bus_w_range49w(0);
	wire_w_lg_w_exp_b_and_w_range72w73w(0) <= wire_w_exp_b_and_w_range72w(0) AND wire_w_exp_b_bus_w_range52w(0);
	wire_w_lg_w_exp_b_and_w_range74w75w(0) <= wire_w_exp_b_and_w_range74w(0) AND wire_w_exp_b_bus_w_range55w(0);
	wire_w_lg_w_exp_b_and_w_range76w77w(0) <= wire_w_exp_b_and_w_range76w(0) AND wire_w_exp_b_bus_w_range58w(0);
	wire_w_lg_w_exp_b_and_w_range78w79w(0) <= wire_w_exp_b_and_w_range78w(0) AND wire_w_exp_b_bus_w_range61w(0);
	wire_w_lg_w_exp_b_and_w_range80w81w(0) <= wire_w_exp_b_and_w_range80w(0) AND wire_w_exp_b_bus_w_range64w(0);
	wire_w_lg_w_exp_bias_and_w_range492w495w(0) <= wire_w_exp_bias_and_w_range492w(0) AND wire_w_exp_bias_bus_w_range494w(0);
	wire_w_lg_w_exp_bias_and_w_range496w498w(0) <= wire_w_exp_bias_and_w_range496w(0) AND wire_w_exp_bias_bus_w_range497w(0);
	wire_w_lg_w_exp_bias_and_w_range499w501w(0) <= wire_w_exp_bias_and_w_range499w(0) AND wire_w_exp_bias_bus_w_range500w(0);
	wire_w_lg_w_exp_bias_and_w_range502w504w(0) <= wire_w_exp_bias_and_w_range502w(0) AND wire_w_exp_bias_bus_w_range503w(0);
	wire_w_lg_w_exp_bias_and_w_range505w507w(0) <= wire_w_exp_bias_and_w_range505w(0) AND wire_w_exp_bias_bus_w_range506w(0);
	wire_w_lg_w_exp_bias_and_w_range508w510w(0) <= wire_w_exp_bias_and_w_range508w(0) AND wire_w_exp_bias_bus_w_range509w(0);
	wire_w_lg_w_exp_bias_and_w_range511w513w(0) <= wire_w_exp_bias_and_w_range511w(0) AND wire_w_exp_bias_bus_w_range512w(0);
	wire_w_lg_w_exp_res_and_w_range680w683w(0) <= wire_w_exp_res_and_w_range680w(0) AND wire_w_exp_res_bus_w_range682w(0);
	wire_w_lg_w_exp_res_and_w_range684w686w(0) <= wire_w_exp_res_and_w_range684w(0) AND wire_w_exp_res_bus_w_range685w(0);
	wire_w_lg_w_exp_res_and_w_range687w689w(0) <= wire_w_exp_res_and_w_range687w(0) AND wire_w_exp_res_bus_w_range688w(0);
	wire_w_lg_w_exp_res_and_w_range690w692w(0) <= wire_w_exp_res_and_w_range690w(0) AND wire_w_exp_res_bus_w_range691w(0);
	wire_w_lg_w_exp_res_and_w_range693w695w(0) <= wire_w_exp_res_and_w_range693w(0) AND wire_w_exp_res_bus_w_range694w(0);
	wire_w_lg_w_exp_res_and_w_range696w698w(0) <= wire_w_exp_res_and_w_range696w(0) AND wire_w_exp_res_bus_w_range697w(0);
	wire_w_lg_w_exp_res_and_w_range699w701w(0) <= wire_w_exp_res_and_w_range699w(0) AND wire_w_exp_res_bus_w_range700w(0);
	wire_w_lg_w_man_a_and_w_range153w155w(0) <= wire_w_man_a_and_w_range153w(0) AND wire_w_man_a_bus_w_range87w(0);
	wire_w_lg_w_man_a_and_w_range174w175w(0) <= wire_w_man_a_and_w_range174w(0) AND wire_w_man_a_bus_w_range117w(0);
	wire_w_lg_w_man_a_and_w_range176w177w(0) <= wire_w_man_a_and_w_range176w(0) AND wire_w_man_a_bus_w_range120w(0);
	wire_w_lg_w_man_a_and_w_range178w179w(0) <= wire_w_man_a_and_w_range178w(0) AND wire_w_man_a_bus_w_range123w(0);
	wire_w_lg_w_man_a_and_w_range180w181w(0) <= wire_w_man_a_and_w_range180w(0) AND wire_w_man_a_bus_w_range126w(0);
	wire_w_lg_w_man_a_and_w_range182w183w(0) <= wire_w_man_a_and_w_range182w(0) AND wire_w_man_a_bus_w_range129w(0);
	wire_w_lg_w_man_a_and_w_range184w185w(0) <= wire_w_man_a_and_w_range184w(0) AND wire_w_man_a_bus_w_range132w(0);
	wire_w_lg_w_man_a_and_w_range186w187w(0) <= wire_w_man_a_and_w_range186w(0) AND wire_w_man_a_bus_w_range135w(0);
	wire_w_lg_w_man_a_and_w_range188w189w(0) <= wire_w_man_a_and_w_range188w(0) AND wire_w_man_a_bus_w_range138w(0);
	wire_w_lg_w_man_a_and_w_range190w191w(0) <= wire_w_man_a_and_w_range190w(0) AND wire_w_man_a_bus_w_range141w(0);
	wire_w_lg_w_man_a_and_w_range192w193w(0) <= wire_w_man_a_and_w_range192w(0) AND wire_w_man_a_bus_w_range144w(0);
	wire_w_lg_w_man_a_and_w_range156w157w(0) <= wire_w_man_a_and_w_range156w(0) AND wire_w_man_a_bus_w_range90w(0);
	wire_w_lg_w_man_a_and_w_range194w195w(0) <= wire_w_man_a_and_w_range194w(0) AND wire_w_man_a_bus_w_range147w(0);
	wire_w_lg_w_man_a_and_w_range196w197w(0) <= wire_w_man_a_and_w_range196w(0) AND wire_w_man_a_bus_w_range150w(0);
	wire_w_lg_w_man_a_and_w_range158w159w(0) <= wire_w_man_a_and_w_range158w(0) AND wire_w_man_a_bus_w_range93w(0);
	wire_w_lg_w_man_a_and_w_range160w161w(0) <= wire_w_man_a_and_w_range160w(0) AND wire_w_man_a_bus_w_range96w(0);
	wire_w_lg_w_man_a_and_w_range162w163w(0) <= wire_w_man_a_and_w_range162w(0) AND wire_w_man_a_bus_w_range99w(0);
	wire_w_lg_w_man_a_and_w_range164w165w(0) <= wire_w_man_a_and_w_range164w(0) AND wire_w_man_a_bus_w_range102w(0);
	wire_w_lg_w_man_a_and_w_range166w167w(0) <= wire_w_man_a_and_w_range166w(0) AND wire_w_man_a_bus_w_range105w(0);
	wire_w_lg_w_man_a_and_w_range168w169w(0) <= wire_w_man_a_and_w_range168w(0) AND wire_w_man_a_bus_w_range108w(0);
	wire_w_lg_w_man_a_and_w_range170w171w(0) <= wire_w_man_a_and_w_range170w(0) AND wire_w_man_a_bus_w_range111w(0);
	wire_w_lg_w_man_a_and_w_range172w173w(0) <= wire_w_man_a_and_w_range172w(0) AND wire_w_man_a_bus_w_range114w(0);
	wire_w_lg_w_man_b_and_w_range269w271w(0) <= wire_w_man_b_and_w_range269w(0) AND wire_w_man_b_bus_w_range203w(0);
	wire_w_lg_w_man_b_and_w_range290w291w(0) <= wire_w_man_b_and_w_range290w(0) AND wire_w_man_b_bus_w_range233w(0);
	wire_w_lg_w_man_b_and_w_range292w293w(0) <= wire_w_man_b_and_w_range292w(0) AND wire_w_man_b_bus_w_range236w(0);
	wire_w_lg_w_man_b_and_w_range294w295w(0) <= wire_w_man_b_and_w_range294w(0) AND wire_w_man_b_bus_w_range239w(0);
	wire_w_lg_w_man_b_and_w_range296w297w(0) <= wire_w_man_b_and_w_range296w(0) AND wire_w_man_b_bus_w_range242w(0);
	wire_w_lg_w_man_b_and_w_range298w299w(0) <= wire_w_man_b_and_w_range298w(0) AND wire_w_man_b_bus_w_range245w(0);
	wire_w_lg_w_man_b_and_w_range300w301w(0) <= wire_w_man_b_and_w_range300w(0) AND wire_w_man_b_bus_w_range248w(0);
	wire_w_lg_w_man_b_and_w_range302w303w(0) <= wire_w_man_b_and_w_range302w(0) AND wire_w_man_b_bus_w_range251w(0);
	wire_w_lg_w_man_b_and_w_range304w305w(0) <= wire_w_man_b_and_w_range304w(0) AND wire_w_man_b_bus_w_range254w(0);
	wire_w_lg_w_man_b_and_w_range306w307w(0) <= wire_w_man_b_and_w_range306w(0) AND wire_w_man_b_bus_w_range257w(0);
	wire_w_lg_w_man_b_and_w_range308w309w(0) <= wire_w_man_b_and_w_range308w(0) AND wire_w_man_b_bus_w_range260w(0);
	wire_w_lg_w_man_b_and_w_range272w273w(0) <= wire_w_man_b_and_w_range272w(0) AND wire_w_man_b_bus_w_range206w(0);
	wire_w_lg_w_man_b_and_w_range310w311w(0) <= wire_w_man_b_and_w_range310w(0) AND wire_w_man_b_bus_w_range263w(0);
	wire_w_lg_w_man_b_and_w_range312w313w(0) <= wire_w_man_b_and_w_range312w(0) AND wire_w_man_b_bus_w_range266w(0);
	wire_w_lg_w_man_b_and_w_range274w275w(0) <= wire_w_man_b_and_w_range274w(0) AND wire_w_man_b_bus_w_range209w(0);
	wire_w_lg_w_man_b_and_w_range276w277w(0) <= wire_w_man_b_and_w_range276w(0) AND wire_w_man_b_bus_w_range212w(0);
	wire_w_lg_w_man_b_and_w_range278w279w(0) <= wire_w_man_b_and_w_range278w(0) AND wire_w_man_b_bus_w_range215w(0);
	wire_w_lg_w_man_b_and_w_range280w281w(0) <= wire_w_man_b_and_w_range280w(0) AND wire_w_man_b_bus_w_range218w(0);
	wire_w_lg_w_man_b_and_w_range282w283w(0) <= wire_w_man_b_and_w_range282w(0) AND wire_w_man_b_bus_w_range221w(0);
	wire_w_lg_w_man_b_and_w_range284w285w(0) <= wire_w_man_b_and_w_range284w(0) AND wire_w_man_b_bus_w_range224w(0);
	wire_w_lg_w_man_b_and_w_range286w287w(0) <= wire_w_man_b_and_w_range286w(0) AND wire_w_man_b_bus_w_range227w(0);
	wire_w_lg_w_man_b_and_w_range288w289w(0) <= wire_w_man_b_and_w_range288w(0) AND wire_w_man_b_bus_w_range230w(0);
	wire_w_lg_w_norm_infi_and_w_range562w565w(0) <= wire_w_norm_infi_and_w_range562w(0) AND wire_w_norm_infi_bus_w_range564w(0);
	wire_w_lg_w_norm_infi_and_w_range566w568w(0) <= wire_w_norm_infi_and_w_range566w(0) AND wire_w_norm_infi_bus_w_range567w(0);
	wire_w_lg_w_norm_infi_and_w_range569w571w(0) <= wire_w_norm_infi_and_w_range569w(0) AND wire_w_norm_infi_bus_w_range570w(0);
	wire_w_lg_w_norm_infi_and_w_range572w574w(0) <= wire_w_norm_infi_and_w_range572w(0) AND wire_w_norm_infi_bus_w_range573w(0);
	wire_w_lg_w_norm_infi_and_w_range575w577w(0) <= wire_w_norm_infi_and_w_range575w(0) AND wire_w_norm_infi_bus_w_range576w(0);
	wire_w_lg_w_norm_infi_and_w_range578w580w(0) <= wire_w_norm_infi_and_w_range578w(0) AND wire_w_norm_infi_bus_w_range579w(0);
	wire_w_lg_w_norm_infi_and_w_range581w583w(0) <= wire_w_norm_infi_and_w_range581w(0) AND wire_w_norm_infi_bus_w_range582w(0);
	wire_w_lg_bias_addition_overf_w521w(0) <= NOT bias_addition_overf_w;
	wire_w_lg_dataa_S0329w(0) <= NOT dataa_S0;
	wire_w_lg_datab_S0339w(0) <= NOT datab_S0;
	wire_w_lg_exp_a_b_w487w(0) <= NOT exp_a_b_w;
	wire_w_lg_exp_a_one_w640w(0) <= NOT exp_a_one_w;
	wire_w_lg_exp_a_or_msb_w325w(0) <= NOT exp_a_or_msb_w;
	wire_w_lg_exp_b_one_w649w(0) <= NOT exp_b_one_w;
	wire_w_lg_exp_b_or_msb_w327w(0) <= NOT exp_b_or_msb_w;
	wire_w_lg_exp_sign_w516w(0) <= NOT exp_sign_w;
	wire_w_lg_guard_bit_dffe1a_w446w(0) <= NOT guard_bit_dffe1a_w;
	wire_w_lg_infi_combi_w779w(0) <= NOT infi_combi_w;
	wire_w_lg_infinite_w800w(0) <= NOT infinite_w;
	wire_w_lg_mux1_exp_s0a475w(0) <= NOT mux1_exp_s0a;
	wire_w_lg_mux1_exp_s1a478w(0) <= NOT mux1_exp_s1a;
	wire_w_lg_mux_zero_non_zero_S0590w(0) <= NOT mux_zero_non_zero_S0;
	wire_w_lg_nan_w780w(0) <= NOT nan_w;
	wire_w_lg_not_exp_res_int2_or_res_w620w(0) <= NOT not_exp_res_int2_or_res_w;
	wire_w_lg_quo_msb_m1_w380w(0) <= NOT quo_msb_m1_w;
	wire_w_lg_rnd_overflow457w(0) <= NOT rnd_overflow;
	wire_w_lg_zero_dataa_w775w(0) <= NOT zero_dataa_w;
	wire_w_lg_zero_w804w(0) <= NOT zero_w;
	wire_w_lg_w_man_res_or_w_range772w773w(0) <= NOT wire_w_man_res_or_w_range772w(0);
	loop102 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_dataa_S0354w355w(i) <= wire_w_lg_dataa_S0354w(i) OR wire_w_lg_w_lg_dataa_S0329w353w(i);
	END GENERATE loop102;
	loop103 : FOR i IN 0 TO 30 GENERATE 
		wire_w_lg_w_lg_datab_S0362w363w(i) <= wire_w_lg_datab_S0362w(i) OR wire_w_lg_w_lg_datab_S0339w361w(i);
	END GENERATE loop103;
	wire_w_lg_w_lg_exp_zero_bus_w587w588w(0) <= wire_w_lg_exp_zero_bus_w587w(0) OR bias_addition_overf_w;
	wire_w_lg_w_lg_man_a_zero_w641w642w(0) <= wire_w_lg_man_a_zero_w641w(0) OR man_a_one_w;
	wire_w_lg_w_lg_man_b_zero_w650w651w(0) <= wire_w_lg_man_b_zero_w650w(0) OR man_b_one_w;
	wire_w_lg_exp_zero_bus_w587w(0) <= exp_zero_bus_w OR signed_N_exp_h_or;
	wire_w_lg_man_a_zero_w641w(0) <= man_a_zero_w OR man_a_non_zero_w;
	wire_w_lg_man_b_zero_w650w(0) <= man_b_zero_w OR man_b_non_zero_w;
	wire_w412w(0) <= sticky_quo_msb_m1_comparator_upper_upper_agb_w OR wire_w411w(0);
	wire_w_lg_w_exp_a_or_w_range3w6w(0) <= wire_w_exp_a_or_w_range3w(0) OR wire_w_exp_a_bus_w_range5w(0);
	wire_w_lg_w_exp_a_or_w_range7w9w(0) <= wire_w_exp_a_or_w_range7w(0) OR wire_w_exp_a_bus_w_range8w(0);
	wire_w_lg_w_exp_a_or_w_range10w12w(0) <= wire_w_exp_a_or_w_range10w(0) OR wire_w_exp_a_bus_w_range11w(0);
	wire_w_lg_w_exp_a_or_w_range13w15w(0) <= wire_w_exp_a_or_w_range13w(0) OR wire_w_exp_a_bus_w_range14w(0);
	wire_w_lg_w_exp_a_or_w_range16w18w(0) <= wire_w_exp_a_or_w_range16w(0) OR wire_w_exp_a_bus_w_range17w(0);
	wire_w_lg_w_exp_a_or_w_range19w21w(0) <= wire_w_exp_a_or_w_range19w(0) OR wire_w_exp_a_bus_w_range20w(0);
	wire_w_lg_w_exp_a_or_w_range22w24w(0) <= wire_w_exp_a_or_w_range22w(0) OR wire_w_exp_a_bus_w_range23w(0);
	wire_w_lg_w_exp_b_or_w_range44w47w(0) <= wire_w_exp_b_or_w_range44w(0) OR wire_w_exp_b_bus_w_range46w(0);
	wire_w_lg_w_exp_b_or_w_range48w50w(0) <= wire_w_exp_b_or_w_range48w(0) OR wire_w_exp_b_bus_w_range49w(0);
	wire_w_lg_w_exp_b_or_w_range51w53w(0) <= wire_w_exp_b_or_w_range51w(0) OR wire_w_exp_b_bus_w_range52w(0);
	wire_w_lg_w_exp_b_or_w_range54w56w(0) <= wire_w_exp_b_or_w_range54w(0) OR wire_w_exp_b_bus_w_range55w(0);
	wire_w_lg_w_exp_b_or_w_range57w59w(0) <= wire_w_exp_b_or_w_range57w(0) OR wire_w_exp_b_bus_w_range58w(0);
	wire_w_lg_w_exp_b_or_w_range60w62w(0) <= wire_w_exp_b_or_w_range60w(0) OR wire_w_exp_b_bus_w_range61w(0);
	wire_w_lg_w_exp_b_or_w_range63w65w(0) <= wire_w_exp_b_or_w_range63w(0) OR wire_w_exp_b_bus_w_range64w(0);
	wire_w_lg_w_exp_higher_or_range531w534w(0) <= wire_w_exp_higher_or_range531w(0) OR wire_w_exp_higher_bit_range533w(0);
	wire_w_lg_w_exp_res_int2_or_w_range596w599w(0) <= wire_w_exp_res_int2_or_w_range596w(0) OR wire_w_exp_res_int2_bus_w_range598w(0);
	wire_w_lg_w_exp_res_int2_or_w_range600w602w(0) <= wire_w_exp_res_int2_or_w_range600w(0) OR wire_w_exp_res_int2_bus_w_range601w(0);
	wire_w_lg_w_exp_res_int2_or_w_range603w605w(0) <= wire_w_exp_res_int2_or_w_range603w(0) OR wire_w_exp_res_int2_bus_w_range604w(0);
	wire_w_lg_w_exp_res_int2_or_w_range606w608w(0) <= wire_w_exp_res_int2_or_w_range606w(0) OR wire_w_exp_res_int2_bus_w_range607w(0);
	wire_w_lg_w_exp_res_int2_or_w_range609w611w(0) <= wire_w_exp_res_int2_or_w_range609w(0) OR wire_w_exp_res_int2_bus_w_range610w(0);
	wire_w_lg_w_exp_res_int2_or_w_range612w614w(0) <= wire_w_exp_res_int2_or_w_range612w(0) OR wire_w_exp_res_int2_bus_w_range613w(0);
	wire_w_lg_w_exp_res_int2_or_w_range615w617w(0) <= wire_w_exp_res_int2_or_w_range615w(0) OR wire_w_exp_res_int2_bus_w_range616w(0);
	wire_w_lg_w_man_a_or_w_range85w88w(0) <= wire_w_man_a_or_w_range85w(0) OR wire_w_man_a_bus_w_range87w(0);
	wire_w_lg_w_man_a_or_w_range116w118w(0) <= wire_w_man_a_or_w_range116w(0) OR wire_w_man_a_bus_w_range117w(0);
	wire_w_lg_w_man_a_or_w_range119w121w(0) <= wire_w_man_a_or_w_range119w(0) OR wire_w_man_a_bus_w_range120w(0);
	wire_w_lg_w_man_a_or_w_range122w124w(0) <= wire_w_man_a_or_w_range122w(0) OR wire_w_man_a_bus_w_range123w(0);
	wire_w_lg_w_man_a_or_w_range125w127w(0) <= wire_w_man_a_or_w_range125w(0) OR wire_w_man_a_bus_w_range126w(0);
	wire_w_lg_w_man_a_or_w_range128w130w(0) <= wire_w_man_a_or_w_range128w(0) OR wire_w_man_a_bus_w_range129w(0);
	wire_w_lg_w_man_a_or_w_range131w133w(0) <= wire_w_man_a_or_w_range131w(0) OR wire_w_man_a_bus_w_range132w(0);
	wire_w_lg_w_man_a_or_w_range134w136w(0) <= wire_w_man_a_or_w_range134w(0) OR wire_w_man_a_bus_w_range135w(0);
	wire_w_lg_w_man_a_or_w_range137w139w(0) <= wire_w_man_a_or_w_range137w(0) OR wire_w_man_a_bus_w_range138w(0);
	wire_w_lg_w_man_a_or_w_range140w142w(0) <= wire_w_man_a_or_w_range140w(0) OR wire_w_man_a_bus_w_range141w(0);
	wire_w_lg_w_man_a_or_w_range143w145w(0) <= wire_w_man_a_or_w_range143w(0) OR wire_w_man_a_bus_w_range144w(0);
	wire_w_lg_w_man_a_or_w_range89w91w(0) <= wire_w_man_a_or_w_range89w(0) OR wire_w_man_a_bus_w_range90w(0);
	wire_w_lg_w_man_a_or_w_range146w148w(0) <= wire_w_man_a_or_w_range146w(0) OR wire_w_man_a_bus_w_range147w(0);
	wire_w_lg_w_man_a_or_w_range149w151w(0) <= wire_w_man_a_or_w_range149w(0) OR wire_w_man_a_bus_w_range150w(0);
	wire_w_lg_w_man_a_or_w_range92w94w(0) <= wire_w_man_a_or_w_range92w(0) OR wire_w_man_a_bus_w_range93w(0);
	wire_w_lg_w_man_a_or_w_range95w97w(0) <= wire_w_man_a_or_w_range95w(0) OR wire_w_man_a_bus_w_range96w(0);
	wire_w_lg_w_man_a_or_w_range98w100w(0) <= wire_w_man_a_or_w_range98w(0) OR wire_w_man_a_bus_w_range99w(0);
	wire_w_lg_w_man_a_or_w_range101w103w(0) <= wire_w_man_a_or_w_range101w(0) OR wire_w_man_a_bus_w_range102w(0);
	wire_w_lg_w_man_a_or_w_range104w106w(0) <= wire_w_man_a_or_w_range104w(0) OR wire_w_man_a_bus_w_range105w(0);
	wire_w_lg_w_man_a_or_w_range107w109w(0) <= wire_w_man_a_or_w_range107w(0) OR wire_w_man_a_bus_w_range108w(0);
	wire_w_lg_w_man_a_or_w_range110w112w(0) <= wire_w_man_a_or_w_range110w(0) OR wire_w_man_a_bus_w_range111w(0);
	wire_w_lg_w_man_a_or_w_range113w115w(0) <= wire_w_man_a_or_w_range113w(0) OR wire_w_man_a_bus_w_range114w(0);
	wire_w_lg_w_man_b_or_w_range201w204w(0) <= wire_w_man_b_or_w_range201w(0) OR wire_w_man_b_bus_w_range203w(0);
	wire_w_lg_w_man_b_or_w_range232w234w(0) <= wire_w_man_b_or_w_range232w(0) OR wire_w_man_b_bus_w_range233w(0);
	wire_w_lg_w_man_b_or_w_range235w237w(0) <= wire_w_man_b_or_w_range235w(0) OR wire_w_man_b_bus_w_range236w(0);
	wire_w_lg_w_man_b_or_w_range238w240w(0) <= wire_w_man_b_or_w_range238w(0) OR wire_w_man_b_bus_w_range239w(0);
	wire_w_lg_w_man_b_or_w_range241w243w(0) <= wire_w_man_b_or_w_range241w(0) OR wire_w_man_b_bus_w_range242w(0);
	wire_w_lg_w_man_b_or_w_range244w246w(0) <= wire_w_man_b_or_w_range244w(0) OR wire_w_man_b_bus_w_range245w(0);
	wire_w_lg_w_man_b_or_w_range247w249w(0) <= wire_w_man_b_or_w_range247w(0) OR wire_w_man_b_bus_w_range248w(0);
	wire_w_lg_w_man_b_or_w_range250w252w(0) <= wire_w_man_b_or_w_range250w(0) OR wire_w_man_b_bus_w_range251w(0);
	wire_w_lg_w_man_b_or_w_range253w255w(0) <= wire_w_man_b_or_w_range253w(0) OR wire_w_man_b_bus_w_range254w(0);
	wire_w_lg_w_man_b_or_w_range256w258w(0) <= wire_w_man_b_or_w_range256w(0) OR wire_w_man_b_bus_w_range257w(0);
	wire_w_lg_w_man_b_or_w_range259w261w(0) <= wire_w_man_b_or_w_range259w(0) OR wire_w_man_b_bus_w_range260w(0);
	wire_w_lg_w_man_b_or_w_range205w207w(0) <= wire_w_man_b_or_w_range205w(0) OR wire_w_man_b_bus_w_range206w(0);
	wire_w_lg_w_man_b_or_w_range262w264w(0) <= wire_w_man_b_or_w_range262w(0) OR wire_w_man_b_bus_w_range263w(0);
	wire_w_lg_w_man_b_or_w_range265w267w(0) <= wire_w_man_b_or_w_range265w(0) OR wire_w_man_b_bus_w_range266w(0);
	wire_w_lg_w_man_b_or_w_range208w210w(0) <= wire_w_man_b_or_w_range208w(0) OR wire_w_man_b_bus_w_range209w(0);
	wire_w_lg_w_man_b_or_w_range211w213w(0) <= wire_w_man_b_or_w_range211w(0) OR wire_w_man_b_bus_w_range212w(0);
	wire_w_lg_w_man_b_or_w_range214w216w(0) <= wire_w_man_b_or_w_range214w(0) OR wire_w_man_b_bus_w_range215w(0);
	wire_w_lg_w_man_b_or_w_range217w219w(0) <= wire_w_man_b_or_w_range217w(0) OR wire_w_man_b_bus_w_range218w(0);
	wire_w_lg_w_man_b_or_w_range220w222w(0) <= wire_w_man_b_or_w_range220w(0) OR wire_w_man_b_bus_w_range221w(0);
	wire_w_lg_w_man_b_or_w_range223w225w(0) <= wire_w_man_b_or_w_range223w(0) OR wire_w_man_b_bus_w_range224w(0);
	wire_w_lg_w_man_b_or_w_range226w228w(0) <= wire_w_man_b_or_w_range226w(0) OR wire_w_man_b_bus_w_range227w(0);
	wire_w_lg_w_man_b_or_w_range229w231w(0) <= wire_w_man_b_or_w_range229w(0) OR wire_w_man_b_bus_w_range230w(0);
	wire_w_lg_w_man_res_or_w_range705w708w(0) <= wire_w_man_res_or_w_range705w(0) OR wire_w_man_res_bus_w_range707w(0);
	wire_w_lg_w_man_res_or_w_range736w738w(0) <= wire_w_man_res_or_w_range736w(0) OR wire_w_man_res_bus_w_range737w(0);
	wire_w_lg_w_man_res_or_w_range739w741w(0) <= wire_w_man_res_or_w_range739w(0) OR wire_w_man_res_bus_w_range740w(0);
	wire_w_lg_w_man_res_or_w_range742w744w(0) <= wire_w_man_res_or_w_range742w(0) OR wire_w_man_res_bus_w_range743w(0);
	wire_w_lg_w_man_res_or_w_range745w747w(0) <= wire_w_man_res_or_w_range745w(0) OR wire_w_man_res_bus_w_range746w(0);
	wire_w_lg_w_man_res_or_w_range748w750w(0) <= wire_w_man_res_or_w_range748w(0) OR wire_w_man_res_bus_w_range749w(0);
	wire_w_lg_w_man_res_or_w_range751w753w(0) <= wire_w_man_res_or_w_range751w(0) OR wire_w_man_res_bus_w_range752w(0);
	wire_w_lg_w_man_res_or_w_range754w756w(0) <= wire_w_man_res_or_w_range754w(0) OR wire_w_man_res_bus_w_range755w(0);
	wire_w_lg_w_man_res_or_w_range757w759w(0) <= wire_w_man_res_or_w_range757w(0) OR wire_w_man_res_bus_w_range758w(0);
	wire_w_lg_w_man_res_or_w_range760w762w(0) <= wire_w_man_res_or_w_range760w(0) OR wire_w_man_res_bus_w_range761w(0);
	wire_w_lg_w_man_res_or_w_range763w765w(0) <= wire_w_man_res_or_w_range763w(0) OR wire_w_man_res_bus_w_range764w(0);
	wire_w_lg_w_man_res_or_w_range709w711w(0) <= wire_w_man_res_or_w_range709w(0) OR wire_w_man_res_bus_w_range710w(0);
	wire_w_lg_w_man_res_or_w_range766w768w(0) <= wire_w_man_res_or_w_range766w(0) OR wire_w_man_res_bus_w_range767w(0);
	wire_w_lg_w_man_res_or_w_range769w771w(0) <= wire_w_man_res_or_w_range769w(0) OR wire_w_man_res_bus_w_range770w(0);
	wire_w_lg_w_man_res_or_w_range712w714w(0) <= wire_w_man_res_or_w_range712w(0) OR wire_w_man_res_bus_w_range713w(0);
	wire_w_lg_w_man_res_or_w_range715w717w(0) <= wire_w_man_res_or_w_range715w(0) OR wire_w_man_res_bus_w_range716w(0);
	wire_w_lg_w_man_res_or_w_range718w720w(0) <= wire_w_man_res_or_w_range718w(0) OR wire_w_man_res_bus_w_range719w(0);
	wire_w_lg_w_man_res_or_w_range721w723w(0) <= wire_w_man_res_or_w_range721w(0) OR wire_w_man_res_bus_w_range722w(0);
	wire_w_lg_w_man_res_or_w_range724w726w(0) <= wire_w_man_res_or_w_range724w(0) OR wire_w_man_res_bus_w_range725w(0);
	wire_w_lg_w_man_res_or_w_range727w729w(0) <= wire_w_man_res_or_w_range727w(0) OR wire_w_man_res_bus_w_range728w(0);
	wire_w_lg_w_man_res_or_w_range730w732w(0) <= wire_w_man_res_or_w_range730w(0) OR wire_w_man_res_bus_w_range731w(0);
	wire_w_lg_w_man_res_or_w_range733w735w(0) <= wire_w_man_res_or_w_range733w(0) OR wire_w_man_res_bus_w_range734w(0);
	wire_w_lg_w_norm_zero_or_w_range537w540w(0) <= wire_w_norm_zero_or_w_range537w(0) OR wire_w_norm_zero_bus_w_range539w(0);
	wire_w_lg_w_norm_zero_or_w_range541w543w(0) <= wire_w_norm_zero_or_w_range541w(0) OR wire_w_norm_zero_bus_w_range542w(0);
	wire_w_lg_w_norm_zero_or_w_range544w546w(0) <= wire_w_norm_zero_or_w_range544w(0) OR wire_w_norm_zero_bus_w_range545w(0);
	wire_w_lg_w_norm_zero_or_w_range547w549w(0) <= wire_w_norm_zero_or_w_range547w(0) OR wire_w_norm_zero_bus_w_range548w(0);
	wire_w_lg_w_norm_zero_or_w_range550w552w(0) <= wire_w_norm_zero_or_w_range550w(0) OR wire_w_norm_zero_bus_w_range551w(0);
	wire_w_lg_w_norm_zero_or_w_range553w555w(0) <= wire_w_norm_zero_or_w_range553w(0) OR wire_w_norm_zero_bus_w_range554w(0);
	wire_w_lg_w_norm_zero_or_w_range556w558w(0) <= wire_w_norm_zero_or_w_range556w(0) OR wire_w_norm_zero_bus_w_range557w(0);
	wire_w_lg_w_sticky_bit_quo_msb_m1_or_range388w391w(0) <= wire_w_sticky_bit_quo_msb_m1_or_range388w(0) OR wire_w_sticky_bit_quo_msb_m1_bit_range390w(0);
	aclr <= '0';
	add_1_dataa_w <= ( checked_quotient_dffe1a_w);
	add_1_datab_w <= (OTHERS => '0');
	add_1_w <= (wire_w_lg_w_lg_w_lg_guard_bit_dffe1a_w446w447w448w(0) OR (guard_bit_dffe1a_w AND round_bit_dffe1a_w));
	add_one_process_w <= wire_altfp_div_csa8_result;
	and_or_dffe1a_w <= and_or_dffe1a;
	and_or_dffe3a_w <= and_or_dffe3a;
	and_or_dffe_w <= and_or_dffe;
	and_or_int_w <= and_or_dffe1a;
	and_or_pipeline_w <= and_or_pipeline27c;
	bias_add_w <= (wire_w_lg_w_lg_exp_a_b_w487w488w OR wire_w_lg_exp_a_b_w486w);
	bias_addition_overf_w <= (wire_add_sub10_overflow OR (wire_w_lg_exp_sign_w516w(0) AND exp_bias_and_res_w));
	bias_addition_w <= wire_add_sub10_result(7 DOWNTO 0);
	bias_value_w <= (((wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w481w482w OR wire_w_lg_w_lg_w_lg_mux1_exp_s1a478w479w480w) OR wire_w_lg_w_lg_mux1_exp_s1a476w477w) OR wire_w_lg_w_lg_mux1_exp_s1a473w474w);
	checked_quotient_dffe1a_w <= checked_quotient_w;
	checked_quotient_w <= (wire_w_lg_quo_msb_m1_w382w OR wire_w_lg_w_lg_quo_msb_m1_w380w381w);
	clk_en <= '1';
	dataa_exp_bus_w <= dataa(30 DOWNTO 23);
	dataa_int <= ( dataa(31) & wire_w_lg_w_lg_dataa_S0354w355w);
	dataa_man_bus_w <= dataa(22 DOWNTO 0);
	dataa_S0 <= (wire_w_lg_exp_a_or_msb_w325w(0) AND man_a_or_msb_w);
	datab_exp_bus_w <= datab(30 DOWNTO 23);
	datab_int <= ( datab(31) & wire_w_lg_w_lg_datab_S0362w363w);
	datab_man_bus_w <= datab(22 DOWNTO 0);
	datab_S0 <= (wire_w_lg_exp_b_or_msb_w327w(0) AND man_b_or_msb_w);
	divider_srt_w <= divider_pipe1a;
	division_by_w <= ((norm_dataa_w AND wire_w_lg_zero_dataa_w775w(0)) AND zero_datab_w);
	division_by_zero <= division_by_zero_port_dffe;
	exp_a_and_msb2_w <= and_or_dffe3a_w(6);
	exp_a_and_msb_w <= exp_a_and_w(7);
	exp_a_and_mux_w <= ((dataa_S0 AND zero_bit_w) OR wire_w_lg_w_lg_dataa_S0329w333w(0));
	exp_a_and_w <= ( wire_w_lg_w_exp_a_and_w_range39w40w & wire_w_lg_w_exp_a_and_w_range37w38w & wire_w_lg_w_exp_a_and_w_range35w36w & wire_w_lg_w_exp_a_and_w_range33w34w & wire_w_lg_w_exp_a_and_w_range31w32w & wire_w_lg_w_exp_a_and_w_range29w30w & wire_w_lg_w_exp_a_and_w_range26w28w & exp_a_bus_w(0));
	exp_a_b_w <= exp_a_b_dffe;
	exp_a_bus_w <= dataa_exp_bus_w;
	exp_a_non_zero_w <= exp_a_or_dffe;
	exp_a_one_w <= exp_a_and_dffe;
	exp_a_or_msb2_w <= and_or_dffe3a_w(7);
	exp_a_or_msb_w <= exp_a_or_w(7);
	exp_a_or_mux_w <= ((dataa_S0 AND zero_bit_w) OR wire_w_lg_w_lg_dataa_S0329w330w(0));
	exp_a_or_w <= ( wire_w_lg_w_exp_a_or_w_range22w24w & wire_w_lg_w_exp_a_or_w_range19w21w & wire_w_lg_w_exp_a_or_w_range16w18w & wire_w_lg_w_exp_a_or_w_range13w15w & wire_w_lg_w_exp_a_or_w_range10w12w & wire_w_lg_w_exp_a_or_w_range7w9w & wire_w_lg_w_exp_a_or_w_range3w6w & exp_a_bus_w(0));
	exp_a_w <= exp_a_dffe;
	exp_a_zero_w <= wire_exp_a_or_dffe_w_lg_q629w(0);
	exp_b_and_msb2_w <= and_or_dffe3a_w(2);
	exp_b_and_msb_w <= exp_b_and_w(7);
	exp_b_and_mux_w <= ((datab_S0 AND zero_bit_w) OR wire_w_lg_w_lg_datab_S0339w343w(0));
	exp_b_and_w <= ( wire_w_lg_w_exp_b_and_w_range80w81w & wire_w_lg_w_exp_b_and_w_range78w79w & wire_w_lg_w_exp_b_and_w_range76w77w & wire_w_lg_w_exp_b_and_w_range74w75w & wire_w_lg_w_exp_b_and_w_range72w73w & wire_w_lg_w_exp_b_and_w_range70w71w & wire_w_lg_w_exp_b_and_w_range67w69w & exp_b_bus_w(0));
	exp_b_bus_w <= datab_exp_bus_w;
	exp_b_non_zero_w <= exp_b_or_dffe;
	exp_b_one_w <= exp_b_and_dffe;
	exp_b_or_msb2_w <= and_or_dffe3a_w(3);
	exp_b_or_msb_w <= exp_b_or_w(7);
	exp_b_or_mux_w <= ((datab_S0 AND zero_bit_w) OR wire_w_lg_w_lg_datab_S0339w340w(0));
	exp_b_or_w <= ( wire_w_lg_w_exp_b_or_w_range63w65w & wire_w_lg_w_exp_b_or_w_range60w62w & wire_w_lg_w_exp_b_or_w_range57w59w & wire_w_lg_w_exp_b_or_w_range54w56w & wire_w_lg_w_exp_b_or_w_range51w53w & wire_w_lg_w_exp_b_or_w_range48w50w & wire_w_lg_w_exp_b_or_w_range44w47w & exp_b_bus_w(0));
	exp_b_w <= exp_b_dffe;
	exp_b_zero_w <= wire_exp_b_or_dffe_w_lg_q632w(0);
	exp_bias_and_res_w <= exp_bias_and_w(7);
	exp_bias_and_w <= ( wire_w_lg_w_exp_bias_and_w_range511w513w & wire_w_lg_w_exp_bias_and_w_range508w510w & wire_w_lg_w_exp_bias_and_w_range505w507w & wire_w_lg_w_exp_bias_and_w_range502w504w & wire_w_lg_w_exp_bias_and_w_range499w501w & wire_w_lg_w_exp_bias_and_w_range496w498w & wire_w_lg_w_exp_bias_and_w_range492w495w & exp_bias_bus_w(0));
	exp_bias_bus_w <= wire_add_sub10_result(7 DOWNTO 0);
	exp_dffe1a_w <= exp_dffe1a;
	exp_dffe2a_w <= exp_dffe2a;
	exp_exc_ones_w <= (OTHERS => '1');
	exp_exc_zeros_w <= (OTHERS => '0');
	exp_higher_bit <= not_bias_addition_w(7 DOWNTO 6);
	exp_higher_or <= ( wire_w_lg_w_exp_higher_or_range531w534w & exp_higher_bit(0));
	exp_infi_bus_w <= norm_infi_and_w(7);
	exp_man_and_or_w <= ( exp_a_or_mux_w & exp_a_and_mux_w & man_a_or_mux_w & man_a_and_mux_w & exp_b_or_mux_w & exp_b_and_mux_w & man_b_or_mux_w & man_b_and_mux_w);
	exp_or_result_w <= (and_or_dffe1a_w(7) OR and_or_dffe1a_w(3));
	exp_pipeline_w <= exp_pipeline26c;
	exp_res_and_w <= ( wire_w_lg_w_exp_res_and_w_range699w701w & wire_w_lg_w_exp_res_and_w_range696w698w & wire_w_lg_w_exp_res_and_w_range693w695w & wire_w_lg_w_exp_res_and_w_range690w692w & wire_w_lg_w_exp_res_and_w_range687w689w & wire_w_lg_w_exp_res_and_w_range684w686w & wire_w_lg_w_exp_res_and_w_range680w683w & exp_res_bus_w(0));
	exp_res_bus_w <= exp_res_w;
	exp_res_int2_bus_w <= exp_res_int2_w;
	exp_res_int2_or_w <= ( wire_w_lg_w_exp_res_int2_or_w_range615w617w & wire_w_lg_w_exp_res_int2_or_w_range612w614w & wire_w_lg_w_exp_res_int2_or_w_range609w611w & wire_w_lg_w_exp_res_int2_or_w_range606w608w & wire_w_lg_w_exp_res_int2_or_w_range603w605w & wire_w_lg_w_exp_res_int2_or_w_range600w602w & wire_w_lg_w_exp_res_int2_or_w_range596w599w & exp_res_int2_bus_w(0));
	exp_res_int2_w <= exp_res_pipe3;
	exp_res_int_w <= ((wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w524w525w OR wire_w_lg_w_lg_w_lg_bias_addition_overf_w521w522w523w) OR wire_w_lg_w_lg_bias_addition_overf_w519w520w);
	exp_res_w <= (wire_w_lg_not_exp_res_int2_or_res_w622w OR wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w621w);
	exp_sign_w <= wire_add_sub10_result(8);
	exp_sub_a_w <= ( "0" & exp_a_w);
	exp_sub_b_w <= ( "0" & exp_b_w);
	exp_sub_w <= wire_add_sub9_result;
	exp_zero_bus_w <= (NOT norm_zero_or_w(7));
	guard_bit_dffe1a_w <= guard_bit_w;
	guard_bit_quo_msb_m1 <= quotient_w(3);
	guard_bit_quo_msb_m2 <= quotient_w(2);
	guard_bit_w <= ((quo_msb_m1_w AND guard_bit_quo_msb_m1) OR wire_w_lg_w_lg_quo_msb_m1_w380w436w(0));
	infi_combi_w <= (((infi_dataa_w AND norm_datab_w) OR (norm_dataa_w AND zero_datab_w)) OR (infi_dataa_w AND zero_datab_w));
	infi_dataa_w <= (exp_a_one_w AND man_a_zero_w);
	infi_datab_w <= (exp_b_one_w AND man_b_zero_w);
	infi_res_w <= ( sign_exc_bit_w & exp_exc_ones_w & man_exc_zeros_w);
	infinite_int_w <= (infi_combi_w OR overflow_int_w);
	infinite_w <= infinite_int_w;
	man_24_zeros_w <= (OTHERS => '0');
	man_a_and_msb2_w <= and_or_dffe3a_w(4);
	man_a_and_msb_w <= man_a_and_w(22);
	man_a_and_mux_w <= ((dataa_S0 AND zero_bit_w) OR wire_w_lg_w_lg_dataa_S0329w337w(0));
	man_a_and_w <= ( wire_w_lg_w_man_a_and_w_range196w197w & wire_w_lg_w_man_a_and_w_range194w195w & wire_w_lg_w_man_a_and_w_range192w193w & wire_w_lg_w_man_a_and_w_range190w191w & wire_w_lg_w_man_a_and_w_range188w189w & wire_w_lg_w_man_a_and_w_range186w187w & wire_w_lg_w_man_a_and_w_range184w185w & wire_w_lg_w_man_a_and_w_range182w183w & wire_w_lg_w_man_a_and_w_range180w181w & wire_w_lg_w_man_a_and_w_range178w179w & wire_w_lg_w_man_a_and_w_range176w177w & wire_w_lg_w_man_a_and_w_range174w175w & wire_w_lg_w_man_a_and_w_range172w173w & wire_w_lg_w_man_a_and_w_range170w171w & wire_w_lg_w_man_a_and_w_range168w169w & wire_w_lg_w_man_a_and_w_range166w167w & wire_w_lg_w_man_a_and_w_range164w165w & wire_w_lg_w_man_a_and_w_range162w163w & wire_w_lg_w_man_a_and_w_range160w161w & wire_w_lg_w_man_a_and_w_range158w159w & wire_w_lg_w_man_a_and_w_range156w157w & wire_w_lg_w_man_a_and_w_range153w155w & man_a_bus_w(0));
	man_a_bus_w <= dataa_man_bus_w;
	man_a_int_w <= man_a_dffe;
	man_a_non_zero_w <= man_a_or_dffe;
	man_a_one_w <= man_a_and_dffe;
	man_a_or_msb2_w <= and_or_dffe3a_w(5);
	man_a_or_msb_w <= man_a_or_w(22);
	man_a_or_mux_w <= ((dataa_S0 AND zero_bit_w) OR wire_w_lg_w_lg_dataa_S0329w335w(0));
	man_a_or_w <= ( wire_w_lg_w_man_a_or_w_range149w151w & wire_w_lg_w_man_a_or_w_range146w148w & wire_w_lg_w_man_a_or_w_range143w145w & wire_w_lg_w_man_a_or_w_range140w142w & wire_w_lg_w_man_a_or_w_range137w139w & wire_w_lg_w_man_a_or_w_range134w136w & wire_w_lg_w_man_a_or_w_range131w133w & wire_w_lg_w_man_a_or_w_range128w130w & wire_w_lg_w_man_a_or_w_range125w127w & wire_w_lg_w_man_a_or_w_range122w124w & wire_w_lg_w_man_a_or_w_range119w121w & wire_w_lg_w_man_a_or_w_range116w118w & wire_w_lg_w_man_a_or_w_range113w115w & wire_w_lg_w_man_a_or_w_range110w112w & wire_w_lg_w_man_a_or_w_range107w109w & wire_w_lg_w_man_a_or_w_range104w106w & wire_w_lg_w_man_a_or_w_range101w103w & wire_w_lg_w_man_a_or_w_range98w100w & wire_w_lg_w_man_a_or_w_range95w97w & wire_w_lg_w_man_a_or_w_range92w94w & wire_w_lg_w_man_a_or_w_range89w91w & wire_w_lg_w_man_a_or_w_range85w88w & man_a_bus_w(0));
	man_a_w <= ( "1" & man_a_int_w);
	man_a_zero_w <= wire_man_a_or_dffe_w_lg_q635w(0);
	man_b_and_msb2_w <= and_or_dffe3a_w(0);
	man_b_and_msb_w <= man_b_and_w(22);
	man_b_and_mux_w <= ((datab_S0 AND zero_bit_w) OR wire_w_lg_w_lg_datab_S0339w347w(0));
	man_b_and_w <= ( wire_w_lg_w_man_b_and_w_range312w313w & wire_w_lg_w_man_b_and_w_range310w311w & wire_w_lg_w_man_b_and_w_range308w309w & wire_w_lg_w_man_b_and_w_range306w307w & wire_w_lg_w_man_b_and_w_range304w305w & wire_w_lg_w_man_b_and_w_range302w303w & wire_w_lg_w_man_b_and_w_range300w301w & wire_w_lg_w_man_b_and_w_range298w299w & wire_w_lg_w_man_b_and_w_range296w297w & wire_w_lg_w_man_b_and_w_range294w295w & wire_w_lg_w_man_b_and_w_range292w293w & wire_w_lg_w_man_b_and_w_range290w291w & wire_w_lg_w_man_b_and_w_range288w289w & wire_w_lg_w_man_b_and_w_range286w287w & wire_w_lg_w_man_b_and_w_range284w285w & wire_w_lg_w_man_b_and_w_range282w283w & wire_w_lg_w_man_b_and_w_range280w281w & wire_w_lg_w_man_b_and_w_range278w279w & wire_w_lg_w_man_b_and_w_range276w277w & wire_w_lg_w_man_b_and_w_range274w275w & wire_w_lg_w_man_b_and_w_range272w273w & wire_w_lg_w_man_b_and_w_range269w271w & man_b_bus_w(0));
	man_b_bus_w <= datab_man_bus_w;
	man_b_int_w <= man_b_dffe;
	man_b_non_zero_w <= man_b_or_dffe;
	man_b_one_w <= man_b_and_dffe;
	man_b_or_msb2_w <= and_or_dffe3a_w(1);
	man_b_or_msb_w <= man_b_or_w(22);
	man_b_or_mux_w <= ((datab_S0 AND zero_bit_w) OR wire_w_lg_w_lg_datab_S0339w345w(0));
	man_b_or_w <= ( wire_w_lg_w_man_b_or_w_range265w267w & wire_w_lg_w_man_b_or_w_range262w264w & wire_w_lg_w_man_b_or_w_range259w261w & wire_w_lg_w_man_b_or_w_range256w258w & wire_w_lg_w_man_b_or_w_range253w255w & wire_w_lg_w_man_b_or_w_range250w252w & wire_w_lg_w_man_b_or_w_range247w249w & wire_w_lg_w_man_b_or_w_range244w246w & wire_w_lg_w_man_b_or_w_range241w243w & wire_w_lg_w_man_b_or_w_range238w240w & wire_w_lg_w_man_b_or_w_range235w237w & wire_w_lg_w_man_b_or_w_range232w234w & wire_w_lg_w_man_b_or_w_range229w231w & wire_w_lg_w_man_b_or_w_range226w228w & wire_w_lg_w_man_b_or_w_range223w225w & wire_w_lg_w_man_b_or_w_range220w222w & wire_w_lg_w_man_b_or_w_range217w219w & wire_w_lg_w_man_b_or_w_range214w216w & wire_w_lg_w_man_b_or_w_range211w213w & wire_w_lg_w_man_b_or_w_range208w210w & wire_w_lg_w_man_b_or_w_range205w207w & wire_w_lg_w_man_b_or_w_range201w204w & man_b_bus_w(0));
	man_b_w <= ( "1" & man_b_int_w);
	man_b_zero_w <= wire_man_b_or_dffe_w_lg_q638w(0);
	man_exc_nan_w <= ( "1" & man_exc_zeros_w(21 DOWNTO 0));
	man_exc_zeros_w <= (OTHERS => '0');
	man_res_bus_w <= man_res_w(22 DOWNTO 0);
	man_res_int2_w <= man_res_pipe3;
	man_res_int_w <= mux_zero_non_zero_w;
	man_res_or_w <= ( wire_w_lg_w_man_res_or_w_range769w771w & wire_w_lg_w_man_res_or_w_range766w768w & wire_w_lg_w_man_res_or_w_range763w765w & wire_w_lg_w_man_res_or_w_range760w762w & wire_w_lg_w_man_res_or_w_range757w759w & wire_w_lg_w_man_res_or_w_range754w756w & wire_w_lg_w_man_res_or_w_range751w753w & wire_w_lg_w_man_res_or_w_range748w750w & wire_w_lg_w_man_res_or_w_range745w747w & wire_w_lg_w_man_res_or_w_range742w744w & wire_w_lg_w_man_res_or_w_range739w741w & wire_w_lg_w_man_res_or_w_range736w738w & wire_w_lg_w_man_res_or_w_range733w735w & wire_w_lg_w_man_res_or_w_range730w732w & wire_w_lg_w_man_res_or_w_range727w729w & wire_w_lg_w_man_res_or_w_range724w726w & wire_w_lg_w_man_res_or_w_range721w723w & wire_w_lg_w_man_res_or_w_range718w720w & wire_w_lg_w_man_res_or_w_range715w717w & wire_w_lg_w_man_res_or_w_range712w714w & wire_w_lg_w_man_res_or_w_range709w711w & wire_w_lg_w_man_res_or_w_range705w708w & man_res_bus_w(0));
	man_res_w <= (wire_w_lg_not_exp_res_int2_or_res_w625w OR wire_w_lg_w_lg_not_exp_res_int2_or_res_w620w624w);
	mux1_exp_s0a <= rnd_add_overf_w;
	mux1_exp_s1a <= implied_bit2a;
	mux_1_res_w <= (wire_w_lg_infinite_w802w OR wire_w_lg_w_lg_infinite_w800w801w);
	mux_2_res_w <= (wire_w_lg_zero_w806w OR wire_w_lg_w_lg_zero_w804w805w);
	mux_3_res_w <= (wire_w_lg_nan_w809w OR wire_w_lg_w_lg_nan_w780w808w);
	mux_zero_non_zero_S0 <= (wire_w_lg_w_lg_exp_zero_bus_w587w588w(0) OR wire_w_lg_exp_infi_bus_w586w(0));
	mux_zero_non_zero_w <= (wire_w_lg_mux_zero_non_zero_S0592w OR wire_w_lg_w_lg_mux_zero_non_zero_S0590w591w);
	nan_dataa_w <= (exp_a_one_w AND (man_a_non_zero_w OR man_a_one_w));
	nan_datab_w <= (exp_b_one_w AND (man_b_non_zero_w OR man_b_one_w));
	nan_res_w <= ( sign_exc_bit_w & exp_exc_ones_w & man_exc_nan_w);
	nan_w <= (((nan_dataa_w OR nan_datab_w) OR (zero_dataa_w AND zero_datab_w)) OR (infi_dataa_w AND infi_datab_w));
	norm_dataa_w <= (wire_w_lg_exp_a_non_zero_w643w(0) AND wire_w_lg_exp_a_one_w640w(0));
	norm_datab_w <= (wire_w_lg_exp_b_non_zero_w652w(0) AND wire_w_lg_exp_b_one_w649w(0));
	norm_infi_and_w <= ( wire_w_lg_w_norm_infi_and_w_range581w583w & wire_w_lg_w_norm_infi_and_w_range578w580w & wire_w_lg_w_norm_infi_and_w_range575w577w & wire_w_lg_w_norm_infi_and_w_range572w574w & wire_w_lg_w_norm_infi_and_w_range569w571w & wire_w_lg_w_norm_infi_and_w_range566w568w & wire_w_lg_w_norm_infi_and_w_range562w565w & norm_infi_bus_w(0));
	norm_infi_bus_w <= bias_addition_w;
	norm_res_int_w <= ( sign_pipe3a & exp_res_w(7 DOWNTO 0) & man_res_w(22 DOWNTO 0));
	norm_zero_bus_w <= bias_addition_w;
	norm_zero_or_w <= ( wire_w_lg_w_norm_zero_or_w_range556w558w & wire_w_lg_w_norm_zero_or_w_range553w555w & wire_w_lg_w_norm_zero_or_w_range550w552w & wire_w_lg_w_norm_zero_or_w_range547w549w & wire_w_lg_w_norm_zero_or_w_range544w546w & wire_w_lg_w_norm_zero_or_w_range541w543w & wire_w_lg_w_norm_zero_or_w_range537w540w & norm_zero_bus_w(0));
	not_bias_addition_w <= (NOT bias_addition_w);
	not_exp_res_int2_or_res_w <= (NOT exp_res_int2_or_w(7));
	overflow_int_w <= ((wire_bias_addition_overf_dffe_w_lg_q781w(0) AND wire_w_lg_infi_combi_w779w(0)) AND (NOT ((norm_dataa_w AND wire_w_lg_zero_dataa_w775w(0)) AND zero_datab_w)));
	overflow_man_w <= ( "1" & "00000000000000000000000");
	overflow_ones_w <= (OTHERS => '1');
	quo_msb_m1_compare_dataa <= ( remainder_srt_w & "00000000000000000000000000000");
	quo_msb_m1_compare_datab <= ( "00000000000000000000000000000" & divider_srt_w);
	quo_msb_m1_compare_w <= ((wire_w412w(0) OR (sticky_quo_msb_m1_comparator_upper_lower_aeb_w AND sticky_quo_msb_m1_comparator_lower_upper_agb_w)) OR (sticky_quo_msb_m1_comparator_lower_upper_aeb_w AND sticky_quo_msb_m1_comparator_lower_lower_ageb_w));
	quo_msb_m1_w <= quotient_w(26);
	quo_msb_m2_compare_dataa <= ( remainder_srt_w & "000000000000000000000000000000");
	quo_msb_m2_compare_datab <= ( "000000000000000000000000000000" & divider_srt_w);
	quo_msb_m2_compare_w <= (sticky_quo_msb_m2_comparator_upper_agb_w OR (sticky_quo_msb_m2_comparator_upper_aeb_w AND sticky_quo_msb_m2_comparator_lower_ageb_w));
	quotient_msb_m1_w <= quotient_w(26 DOWNTO 3);
	quotient_msb_m2_w <= quotient_w(25 DOWNTO 2);
	quotient_w <= quotient_pipe1a;
	remainder_srt_w <= remainder_pipe1a;
	res_rnded_man_w <= rnded_man_pipe2a;
	result <= result_output_dffe;
	rnd_add_overf_w <= rnd_overflow_dffe;
	rnd_overflow <= wire_altfp_div_csa8_cout;
	rnded_man_w <= (wire_w_lg_rnd_overflow459w OR wire_w_lg_w_lg_rnd_overflow457w458w);
	round_bit_dffe1a_w <= round_bit_w;
	round_bit_quo_msb_m1 <= quotient_w(2);
	round_bit_quo_msb_m2 <= quotient_w(1);
	round_bit_w <= ((quo_msb_m1_w AND round_bit_quo_msb_m1) OR wire_w_lg_w_lg_quo_msb_m1_w380w439w(0));
	sign_a_w <= sign_a_dffe;
	sign_b_w <= sign_b_dffe;
	sign_div <= (sign_a_w XOR sign_b_w);
	sign_div_pipeline_w <= sign_div_pipeline27c;
	sign_exc_bit_w <= sign_pipe3a;
	signed_N_exp_h_or <= (exp_sign_w AND exp_higher_or(1));
	sticky_bit_dffe1a_w <= sticky_bit_w;
	sticky_bit_quo_msb_m1 <= (quo_msb_m1_compare_w OR sticky_bit_quo_msb_m1_or(1));
	sticky_bit_quo_msb_m1_bit <= sticky_bit_quo_msb_m1_tmp;
	sticky_bit_quo_msb_m1_or <= ( wire_w_lg_w_sticky_bit_quo_msb_m1_or_range388w391w & sticky_bit_quo_msb_m1_bit(0));
	sticky_bit_quo_msb_m1_tmp <= quotient_w(1 DOWNTO 0);
	sticky_bit_quo_msb_m2 <= (quo_msb_m2_compare_w OR sticky_bit_quo_msb_m2_or(0));
	sticky_bit_quo_msb_m2_bit <= sticky_bit_quo_msb_m2_tmp;
	sticky_bit_quo_msb_m2_or(0) <= ( sticky_bit_quo_msb_m2_bit(0));
	sticky_bit_quo_msb_m2_tmp(0) <= quotient_w(0);
	sticky_bit_w <= ((quo_msb_m1_w AND sticky_bit_quo_msb_m1) OR wire_w_lg_w_lg_quo_msb_m1_w380w442w(0));
	sticky_quo_msb_m1_comparator_lower_lower_ageb_w <= wire_cmpr5_ageb;
	sticky_quo_msb_m1_comparator_lower_upper_aeb_w <= wire_cmpr4_aeb;
	sticky_quo_msb_m1_comparator_lower_upper_agb_w <= wire_cmpr4_agb;
	sticky_quo_msb_m1_comparator_upper_lower_aeb_w <= wire_cmpr3_aeb;
	sticky_quo_msb_m1_comparator_upper_lower_agb_w <= wire_cmpr3_agb;
	sticky_quo_msb_m1_comparator_upper_upper_aeb_w <= wire_cmpr2_aeb;
	sticky_quo_msb_m1_comparator_upper_upper_agb_w <= wire_cmpr2_agb;
	sticky_quo_msb_m2_comparator_lower_ageb_w <= wire_cmpr7_ageb;
	sticky_quo_msb_m2_comparator_upper_aeb_w <= wire_cmpr6_aeb;
	sticky_quo_msb_m2_comparator_upper_agb_w <= wire_cmpr6_agb;
	underflow_zeros_w <= (OTHERS => '0');
	value_add_1_w <= "010000000";
	value_minus_1_w <= "001111110";
	value_normal_w <= "001111111";
	value_zero_w <= (OTHERS => '0');
	zero_bit_23_w <= (OTHERS => '0');
	zero_bit_31_w <= (OTHERS => '0');
	zero_bit_8_w <= (OTHERS => '0');
	zero_bit_w <= '0';
	zero_dataa_w <= (exp_a_zero_w AND man_a_zero_w);
	zero_datab_w <= (exp_b_zero_w AND man_b_zero_w);
	zero_res_w <= ( sign_exc_bit_w & exp_exc_zeros_w & man_exc_zeros_w);
	zero_w <= (((zero_dataa_w AND norm_datab_w) OR (norm_dataa_w AND infi_datab_w)) OR (zero_dataa_w AND infi_datab_w));
	wire_w_dataa_range352w <= dataa(30 DOWNTO 0);
	wire_w_dataa_int_range366w <= dataa_int(22 DOWNTO 0);
	wire_w_dataa_int_range365w <= dataa_int(30 DOWNTO 23);
	wire_w_datab_range360w <= datab(30 DOWNTO 0);
	wire_w_datab_int_range368w <= datab_int(22 DOWNTO 0);
	wire_w_datab_int_range367w <= datab_int(30 DOWNTO 23);
	wire_w_exp_a_and_w_range26w(0) <= exp_a_and_w(0);
	wire_w_exp_a_and_w_range29w(0) <= exp_a_and_w(1);
	wire_w_exp_a_and_w_range31w(0) <= exp_a_and_w(2);
	wire_w_exp_a_and_w_range33w(0) <= exp_a_and_w(3);
	wire_w_exp_a_and_w_range35w(0) <= exp_a_and_w(4);
	wire_w_exp_a_and_w_range37w(0) <= exp_a_and_w(5);
	wire_w_exp_a_and_w_range39w(0) <= exp_a_and_w(6);
	wire_w_exp_a_bus_w_range5w(0) <= exp_a_bus_w(1);
	wire_w_exp_a_bus_w_range8w(0) <= exp_a_bus_w(2);
	wire_w_exp_a_bus_w_range11w(0) <= exp_a_bus_w(3);
	wire_w_exp_a_bus_w_range14w(0) <= exp_a_bus_w(4);
	wire_w_exp_a_bus_w_range17w(0) <= exp_a_bus_w(5);
	wire_w_exp_a_bus_w_range20w(0) <= exp_a_bus_w(6);
	wire_w_exp_a_bus_w_range23w(0) <= exp_a_bus_w(7);
	wire_w_exp_a_or_w_range3w(0) <= exp_a_or_w(0);
	wire_w_exp_a_or_w_range7w(0) <= exp_a_or_w(1);
	wire_w_exp_a_or_w_range10w(0) <= exp_a_or_w(2);
	wire_w_exp_a_or_w_range13w(0) <= exp_a_or_w(3);
	wire_w_exp_a_or_w_range16w(0) <= exp_a_or_w(4);
	wire_w_exp_a_or_w_range19w(0) <= exp_a_or_w(5);
	wire_w_exp_a_or_w_range22w(0) <= exp_a_or_w(6);
	wire_w_exp_b_and_w_range67w(0) <= exp_b_and_w(0);
	wire_w_exp_b_and_w_range70w(0) <= exp_b_and_w(1);
	wire_w_exp_b_and_w_range72w(0) <= exp_b_and_w(2);
	wire_w_exp_b_and_w_range74w(0) <= exp_b_and_w(3);
	wire_w_exp_b_and_w_range76w(0) <= exp_b_and_w(4);
	wire_w_exp_b_and_w_range78w(0) <= exp_b_and_w(5);
	wire_w_exp_b_and_w_range80w(0) <= exp_b_and_w(6);
	wire_w_exp_b_bus_w_range46w(0) <= exp_b_bus_w(1);
	wire_w_exp_b_bus_w_range49w(0) <= exp_b_bus_w(2);
	wire_w_exp_b_bus_w_range52w(0) <= exp_b_bus_w(3);
	wire_w_exp_b_bus_w_range55w(0) <= exp_b_bus_w(4);
	wire_w_exp_b_bus_w_range58w(0) <= exp_b_bus_w(5);
	wire_w_exp_b_bus_w_range61w(0) <= exp_b_bus_w(6);
	wire_w_exp_b_bus_w_range64w(0) <= exp_b_bus_w(7);
	wire_w_exp_b_or_w_range44w(0) <= exp_b_or_w(0);
	wire_w_exp_b_or_w_range48w(0) <= exp_b_or_w(1);
	wire_w_exp_b_or_w_range51w(0) <= exp_b_or_w(2);
	wire_w_exp_b_or_w_range54w(0) <= exp_b_or_w(3);
	wire_w_exp_b_or_w_range57w(0) <= exp_b_or_w(4);
	wire_w_exp_b_or_w_range60w(0) <= exp_b_or_w(5);
	wire_w_exp_b_or_w_range63w(0) <= exp_b_or_w(6);
	wire_w_exp_bias_and_w_range492w(0) <= exp_bias_and_w(0);
	wire_w_exp_bias_and_w_range496w(0) <= exp_bias_and_w(1);
	wire_w_exp_bias_and_w_range499w(0) <= exp_bias_and_w(2);
	wire_w_exp_bias_and_w_range502w(0) <= exp_bias_and_w(3);
	wire_w_exp_bias_and_w_range505w(0) <= exp_bias_and_w(4);
	wire_w_exp_bias_and_w_range508w(0) <= exp_bias_and_w(5);
	wire_w_exp_bias_and_w_range511w(0) <= exp_bias_and_w(6);
	wire_w_exp_bias_bus_w_range494w(0) <= exp_bias_bus_w(1);
	wire_w_exp_bias_bus_w_range497w(0) <= exp_bias_bus_w(2);
	wire_w_exp_bias_bus_w_range500w(0) <= exp_bias_bus_w(3);
	wire_w_exp_bias_bus_w_range503w(0) <= exp_bias_bus_w(4);
	wire_w_exp_bias_bus_w_range506w(0) <= exp_bias_bus_w(5);
	wire_w_exp_bias_bus_w_range509w(0) <= exp_bias_bus_w(6);
	wire_w_exp_bias_bus_w_range512w(0) <= exp_bias_bus_w(7);
	wire_w_exp_higher_bit_range533w(0) <= exp_higher_bit(1);
	wire_w_exp_higher_or_range531w(0) <= exp_higher_or(0);
	wire_w_exp_res_and_w_range680w(0) <= exp_res_and_w(0);
	wire_w_exp_res_and_w_range684w(0) <= exp_res_and_w(1);
	wire_w_exp_res_and_w_range687w(0) <= exp_res_and_w(2);
	wire_w_exp_res_and_w_range690w(0) <= exp_res_and_w(3);
	wire_w_exp_res_and_w_range693w(0) <= exp_res_and_w(4);
	wire_w_exp_res_and_w_range696w(0) <= exp_res_and_w(5);
	wire_w_exp_res_and_w_range699w(0) <= exp_res_and_w(6);
	wire_w_exp_res_and_w_range702w(0) <= exp_res_and_w(7);
	wire_w_exp_res_bus_w_range682w(0) <= exp_res_bus_w(1);
	wire_w_exp_res_bus_w_range685w(0) <= exp_res_bus_w(2);
	wire_w_exp_res_bus_w_range688w(0) <= exp_res_bus_w(3);
	wire_w_exp_res_bus_w_range691w(0) <= exp_res_bus_w(4);
	wire_w_exp_res_bus_w_range694w(0) <= exp_res_bus_w(5);
	wire_w_exp_res_bus_w_range697w(0) <= exp_res_bus_w(6);
	wire_w_exp_res_bus_w_range700w(0) <= exp_res_bus_w(7);
	wire_w_exp_res_int2_bus_w_range598w(0) <= exp_res_int2_bus_w(1);
	wire_w_exp_res_int2_bus_w_range601w(0) <= exp_res_int2_bus_w(2);
	wire_w_exp_res_int2_bus_w_range604w(0) <= exp_res_int2_bus_w(3);
	wire_w_exp_res_int2_bus_w_range607w(0) <= exp_res_int2_bus_w(4);
	wire_w_exp_res_int2_bus_w_range610w(0) <= exp_res_int2_bus_w(5);
	wire_w_exp_res_int2_bus_w_range613w(0) <= exp_res_int2_bus_w(6);
	wire_w_exp_res_int2_bus_w_range616w(0) <= exp_res_int2_bus_w(7);
	wire_w_exp_res_int2_or_w_range596w(0) <= exp_res_int2_or_w(0);
	wire_w_exp_res_int2_or_w_range600w(0) <= exp_res_int2_or_w(1);
	wire_w_exp_res_int2_or_w_range603w(0) <= exp_res_int2_or_w(2);
	wire_w_exp_res_int2_or_w_range606w(0) <= exp_res_int2_or_w(3);
	wire_w_exp_res_int2_or_w_range609w(0) <= exp_res_int2_or_w(4);
	wire_w_exp_res_int2_or_w_range612w(0) <= exp_res_int2_or_w(5);
	wire_w_exp_res_int2_or_w_range615w(0) <= exp_res_int2_or_w(6);
	wire_w_man_a_and_w_range153w(0) <= man_a_and_w(0);
	wire_w_man_a_and_w_range174w(0) <= man_a_and_w(10);
	wire_w_man_a_and_w_range176w(0) <= man_a_and_w(11);
	wire_w_man_a_and_w_range178w(0) <= man_a_and_w(12);
	wire_w_man_a_and_w_range180w(0) <= man_a_and_w(13);
	wire_w_man_a_and_w_range182w(0) <= man_a_and_w(14);
	wire_w_man_a_and_w_range184w(0) <= man_a_and_w(15);
	wire_w_man_a_and_w_range186w(0) <= man_a_and_w(16);
	wire_w_man_a_and_w_range188w(0) <= man_a_and_w(17);
	wire_w_man_a_and_w_range190w(0) <= man_a_and_w(18);
	wire_w_man_a_and_w_range192w(0) <= man_a_and_w(19);
	wire_w_man_a_and_w_range156w(0) <= man_a_and_w(1);
	wire_w_man_a_and_w_range194w(0) <= man_a_and_w(20);
	wire_w_man_a_and_w_range196w(0) <= man_a_and_w(21);
	wire_w_man_a_and_w_range158w(0) <= man_a_and_w(2);
	wire_w_man_a_and_w_range160w(0) <= man_a_and_w(3);
	wire_w_man_a_and_w_range162w(0) <= man_a_and_w(4);
	wire_w_man_a_and_w_range164w(0) <= man_a_and_w(5);
	wire_w_man_a_and_w_range166w(0) <= man_a_and_w(6);
	wire_w_man_a_and_w_range168w(0) <= man_a_and_w(7);
	wire_w_man_a_and_w_range170w(0) <= man_a_and_w(8);
	wire_w_man_a_and_w_range172w(0) <= man_a_and_w(9);
	wire_w_man_a_bus_w_range114w(0) <= man_a_bus_w(10);
	wire_w_man_a_bus_w_range117w(0) <= man_a_bus_w(11);
	wire_w_man_a_bus_w_range120w(0) <= man_a_bus_w(12);
	wire_w_man_a_bus_w_range123w(0) <= man_a_bus_w(13);
	wire_w_man_a_bus_w_range126w(0) <= man_a_bus_w(14);
	wire_w_man_a_bus_w_range129w(0) <= man_a_bus_w(15);
	wire_w_man_a_bus_w_range132w(0) <= man_a_bus_w(16);
	wire_w_man_a_bus_w_range135w(0) <= man_a_bus_w(17);
	wire_w_man_a_bus_w_range138w(0) <= man_a_bus_w(18);
	wire_w_man_a_bus_w_range141w(0) <= man_a_bus_w(19);
	wire_w_man_a_bus_w_range87w(0) <= man_a_bus_w(1);
	wire_w_man_a_bus_w_range144w(0) <= man_a_bus_w(20);
	wire_w_man_a_bus_w_range147w(0) <= man_a_bus_w(21);
	wire_w_man_a_bus_w_range150w(0) <= man_a_bus_w(22);
	wire_w_man_a_bus_w_range90w(0) <= man_a_bus_w(2);
	wire_w_man_a_bus_w_range93w(0) <= man_a_bus_w(3);
	wire_w_man_a_bus_w_range96w(0) <= man_a_bus_w(4);
	wire_w_man_a_bus_w_range99w(0) <= man_a_bus_w(5);
	wire_w_man_a_bus_w_range102w(0) <= man_a_bus_w(6);
	wire_w_man_a_bus_w_range105w(0) <= man_a_bus_w(7);
	wire_w_man_a_bus_w_range108w(0) <= man_a_bus_w(8);
	wire_w_man_a_bus_w_range111w(0) <= man_a_bus_w(9);
	wire_w_man_a_or_w_range85w(0) <= man_a_or_w(0);
	wire_w_man_a_or_w_range116w(0) <= man_a_or_w(10);
	wire_w_man_a_or_w_range119w(0) <= man_a_or_w(11);
	wire_w_man_a_or_w_range122w(0) <= man_a_or_w(12);
	wire_w_man_a_or_w_range125w(0) <= man_a_or_w(13);
	wire_w_man_a_or_w_range128w(0) <= man_a_or_w(14);
	wire_w_man_a_or_w_range131w(0) <= man_a_or_w(15);
	wire_w_man_a_or_w_range134w(0) <= man_a_or_w(16);
	wire_w_man_a_or_w_range137w(0) <= man_a_or_w(17);
	wire_w_man_a_or_w_range140w(0) <= man_a_or_w(18);
	wire_w_man_a_or_w_range143w(0) <= man_a_or_w(19);
	wire_w_man_a_or_w_range89w(0) <= man_a_or_w(1);
	wire_w_man_a_or_w_range146w(0) <= man_a_or_w(20);
	wire_w_man_a_or_w_range149w(0) <= man_a_or_w(21);
	wire_w_man_a_or_w_range92w(0) <= man_a_or_w(2);
	wire_w_man_a_or_w_range95w(0) <= man_a_or_w(3);
	wire_w_man_a_or_w_range98w(0) <= man_a_or_w(4);
	wire_w_man_a_or_w_range101w(0) <= man_a_or_w(5);
	wire_w_man_a_or_w_range104w(0) <= man_a_or_w(6);
	wire_w_man_a_or_w_range107w(0) <= man_a_or_w(7);
	wire_w_man_a_or_w_range110w(0) <= man_a_or_w(8);
	wire_w_man_a_or_w_range113w(0) <= man_a_or_w(9);
	wire_w_man_b_and_w_range269w(0) <= man_b_and_w(0);
	wire_w_man_b_and_w_range290w(0) <= man_b_and_w(10);
	wire_w_man_b_and_w_range292w(0) <= man_b_and_w(11);
	wire_w_man_b_and_w_range294w(0) <= man_b_and_w(12);
	wire_w_man_b_and_w_range296w(0) <= man_b_and_w(13);
	wire_w_man_b_and_w_range298w(0) <= man_b_and_w(14);
	wire_w_man_b_and_w_range300w(0) <= man_b_and_w(15);
	wire_w_man_b_and_w_range302w(0) <= man_b_and_w(16);
	wire_w_man_b_and_w_range304w(0) <= man_b_and_w(17);
	wire_w_man_b_and_w_range306w(0) <= man_b_and_w(18);
	wire_w_man_b_and_w_range308w(0) <= man_b_and_w(19);
	wire_w_man_b_and_w_range272w(0) <= man_b_and_w(1);
	wire_w_man_b_and_w_range310w(0) <= man_b_and_w(20);
	wire_w_man_b_and_w_range312w(0) <= man_b_and_w(21);
	wire_w_man_b_and_w_range274w(0) <= man_b_and_w(2);
	wire_w_man_b_and_w_range276w(0) <= man_b_and_w(3);
	wire_w_man_b_and_w_range278w(0) <= man_b_and_w(4);
	wire_w_man_b_and_w_range280w(0) <= man_b_and_w(5);
	wire_w_man_b_and_w_range282w(0) <= man_b_and_w(6);
	wire_w_man_b_and_w_range284w(0) <= man_b_and_w(7);
	wire_w_man_b_and_w_range286w(0) <= man_b_and_w(8);
	wire_w_man_b_and_w_range288w(0) <= man_b_and_w(9);
	wire_w_man_b_bus_w_range230w(0) <= man_b_bus_w(10);
	wire_w_man_b_bus_w_range233w(0) <= man_b_bus_w(11);
	wire_w_man_b_bus_w_range236w(0) <= man_b_bus_w(12);
	wire_w_man_b_bus_w_range239w(0) <= man_b_bus_w(13);
	wire_w_man_b_bus_w_range242w(0) <= man_b_bus_w(14);
	wire_w_man_b_bus_w_range245w(0) <= man_b_bus_w(15);
	wire_w_man_b_bus_w_range248w(0) <= man_b_bus_w(16);
	wire_w_man_b_bus_w_range251w(0) <= man_b_bus_w(17);
	wire_w_man_b_bus_w_range254w(0) <= man_b_bus_w(18);
	wire_w_man_b_bus_w_range257w(0) <= man_b_bus_w(19);
	wire_w_man_b_bus_w_range203w(0) <= man_b_bus_w(1);
	wire_w_man_b_bus_w_range260w(0) <= man_b_bus_w(20);
	wire_w_man_b_bus_w_range263w(0) <= man_b_bus_w(21);
	wire_w_man_b_bus_w_range266w(0) <= man_b_bus_w(22);
	wire_w_man_b_bus_w_range206w(0) <= man_b_bus_w(2);
	wire_w_man_b_bus_w_range209w(0) <= man_b_bus_w(3);
	wire_w_man_b_bus_w_range212w(0) <= man_b_bus_w(4);
	wire_w_man_b_bus_w_range215w(0) <= man_b_bus_w(5);
	wire_w_man_b_bus_w_range218w(0) <= man_b_bus_w(6);
	wire_w_man_b_bus_w_range221w(0) <= man_b_bus_w(7);
	wire_w_man_b_bus_w_range224w(0) <= man_b_bus_w(8);
	wire_w_man_b_bus_w_range227w(0) <= man_b_bus_w(9);
	wire_w_man_b_or_w_range201w(0) <= man_b_or_w(0);
	wire_w_man_b_or_w_range232w(0) <= man_b_or_w(10);
	wire_w_man_b_or_w_range235w(0) <= man_b_or_w(11);
	wire_w_man_b_or_w_range238w(0) <= man_b_or_w(12);
	wire_w_man_b_or_w_range241w(0) <= man_b_or_w(13);
	wire_w_man_b_or_w_range244w(0) <= man_b_or_w(14);
	wire_w_man_b_or_w_range247w(0) <= man_b_or_w(15);
	wire_w_man_b_or_w_range250w(0) <= man_b_or_w(16);
	wire_w_man_b_or_w_range253w(0) <= man_b_or_w(17);
	wire_w_man_b_or_w_range256w(0) <= man_b_or_w(18);
	wire_w_man_b_or_w_range259w(0) <= man_b_or_w(19);
	wire_w_man_b_or_w_range205w(0) <= man_b_or_w(1);
	wire_w_man_b_or_w_range262w(0) <= man_b_or_w(20);
	wire_w_man_b_or_w_range265w(0) <= man_b_or_w(21);
	wire_w_man_b_or_w_range208w(0) <= man_b_or_w(2);
	wire_w_man_b_or_w_range211w(0) <= man_b_or_w(3);
	wire_w_man_b_or_w_range214w(0) <= man_b_or_w(4);
	wire_w_man_b_or_w_range217w(0) <= man_b_or_w(5);
	wire_w_man_b_or_w_range220w(0) <= man_b_or_w(6);
	wire_w_man_b_or_w_range223w(0) <= man_b_or_w(7);
	wire_w_man_b_or_w_range226w(0) <= man_b_or_w(8);
	wire_w_man_b_or_w_range229w(0) <= man_b_or_w(9);
	wire_w_man_res_bus_w_range734w(0) <= man_res_bus_w(10);
	wire_w_man_res_bus_w_range737w(0) <= man_res_bus_w(11);
	wire_w_man_res_bus_w_range740w(0) <= man_res_bus_w(12);
	wire_w_man_res_bus_w_range743w(0) <= man_res_bus_w(13);
	wire_w_man_res_bus_w_range746w(0) <= man_res_bus_w(14);
	wire_w_man_res_bus_w_range749w(0) <= man_res_bus_w(15);
	wire_w_man_res_bus_w_range752w(0) <= man_res_bus_w(16);
	wire_w_man_res_bus_w_range755w(0) <= man_res_bus_w(17);
	wire_w_man_res_bus_w_range758w(0) <= man_res_bus_w(18);
	wire_w_man_res_bus_w_range761w(0) <= man_res_bus_w(19);
	wire_w_man_res_bus_w_range707w(0) <= man_res_bus_w(1);
	wire_w_man_res_bus_w_range764w(0) <= man_res_bus_w(20);
	wire_w_man_res_bus_w_range767w(0) <= man_res_bus_w(21);
	wire_w_man_res_bus_w_range770w(0) <= man_res_bus_w(22);
	wire_w_man_res_bus_w_range710w(0) <= man_res_bus_w(2);
	wire_w_man_res_bus_w_range713w(0) <= man_res_bus_w(3);
	wire_w_man_res_bus_w_range716w(0) <= man_res_bus_w(4);
	wire_w_man_res_bus_w_range719w(0) <= man_res_bus_w(5);
	wire_w_man_res_bus_w_range722w(0) <= man_res_bus_w(6);
	wire_w_man_res_bus_w_range725w(0) <= man_res_bus_w(7);
	wire_w_man_res_bus_w_range728w(0) <= man_res_bus_w(8);
	wire_w_man_res_bus_w_range731w(0) <= man_res_bus_w(9);
	wire_w_man_res_or_w_range705w(0) <= man_res_or_w(0);
	wire_w_man_res_or_w_range736w(0) <= man_res_or_w(10);
	wire_w_man_res_or_w_range739w(0) <= man_res_or_w(11);
	wire_w_man_res_or_w_range742w(0) <= man_res_or_w(12);
	wire_w_man_res_or_w_range745w(0) <= man_res_or_w(13);
	wire_w_man_res_or_w_range748w(0) <= man_res_or_w(14);
	wire_w_man_res_or_w_range751w(0) <= man_res_or_w(15);
	wire_w_man_res_or_w_range754w(0) <= man_res_or_w(16);
	wire_w_man_res_or_w_range757w(0) <= man_res_or_w(17);
	wire_w_man_res_or_w_range760w(0) <= man_res_or_w(18);
	wire_w_man_res_or_w_range763w(0) <= man_res_or_w(19);
	wire_w_man_res_or_w_range709w(0) <= man_res_or_w(1);
	wire_w_man_res_or_w_range766w(0) <= man_res_or_w(20);
	wire_w_man_res_or_w_range769w(0) <= man_res_or_w(21);
	wire_w_man_res_or_w_range772w(0) <= man_res_or_w(22);
	wire_w_man_res_or_w_range712w(0) <= man_res_or_w(2);
	wire_w_man_res_or_w_range715w(0) <= man_res_or_w(3);
	wire_w_man_res_or_w_range718w(0) <= man_res_or_w(4);
	wire_w_man_res_or_w_range721w(0) <= man_res_or_w(5);
	wire_w_man_res_or_w_range724w(0) <= man_res_or_w(6);
	wire_w_man_res_or_w_range727w(0) <= man_res_or_w(7);
	wire_w_man_res_or_w_range730w(0) <= man_res_or_w(8);
	wire_w_man_res_or_w_range733w(0) <= man_res_or_w(9);
	wire_w_norm_infi_and_w_range562w(0) <= norm_infi_and_w(0);
	wire_w_norm_infi_and_w_range566w(0) <= norm_infi_and_w(1);
	wire_w_norm_infi_and_w_range569w(0) <= norm_infi_and_w(2);
	wire_w_norm_infi_and_w_range572w(0) <= norm_infi_and_w(3);
	wire_w_norm_infi_and_w_range575w(0) <= norm_infi_and_w(4);
	wire_w_norm_infi_and_w_range578w(0) <= norm_infi_and_w(5);
	wire_w_norm_infi_and_w_range581w(0) <= norm_infi_and_w(6);
	wire_w_norm_infi_bus_w_range564w(0) <= norm_infi_bus_w(1);
	wire_w_norm_infi_bus_w_range567w(0) <= norm_infi_bus_w(2);
	wire_w_norm_infi_bus_w_range570w(0) <= norm_infi_bus_w(3);
	wire_w_norm_infi_bus_w_range573w(0) <= norm_infi_bus_w(4);
	wire_w_norm_infi_bus_w_range576w(0) <= norm_infi_bus_w(5);
	wire_w_norm_infi_bus_w_range579w(0) <= norm_infi_bus_w(6);
	wire_w_norm_infi_bus_w_range582w(0) <= norm_infi_bus_w(7);
	wire_w_norm_zero_bus_w_range539w(0) <= norm_zero_bus_w(1);
	wire_w_norm_zero_bus_w_range542w(0) <= norm_zero_bus_w(2);
	wire_w_norm_zero_bus_w_range545w(0) <= norm_zero_bus_w(3);
	wire_w_norm_zero_bus_w_range548w(0) <= norm_zero_bus_w(4);
	wire_w_norm_zero_bus_w_range551w(0) <= norm_zero_bus_w(5);
	wire_w_norm_zero_bus_w_range554w(0) <= norm_zero_bus_w(6);
	wire_w_norm_zero_bus_w_range557w(0) <= norm_zero_bus_w(7);
	wire_w_norm_zero_or_w_range537w(0) <= norm_zero_or_w(0);
	wire_w_norm_zero_or_w_range541w(0) <= norm_zero_or_w(1);
	wire_w_norm_zero_or_w_range544w(0) <= norm_zero_or_w(2);
	wire_w_norm_zero_or_w_range547w(0) <= norm_zero_or_w(3);
	wire_w_norm_zero_or_w_range550w(0) <= norm_zero_or_w(4);
	wire_w_norm_zero_or_w_range553w(0) <= norm_zero_or_w(5);
	wire_w_norm_zero_or_w_range556w(0) <= norm_zero_or_w(6);
	wire_w_sticky_bit_quo_msb_m1_bit_range390w(0) <= sticky_bit_quo_msb_m1_bit(1);
	wire_w_sticky_bit_quo_msb_m1_or_range388w(0) <= sticky_bit_quo_msb_m1_or(0);
	altfp_div_csa8 :  Float_32_Div_altfp_div_csa_gvc
	  PORT MAP ( 
		cin => add_1_w,
		cout => wire_altfp_div_csa8_cout,
		dataa => add_1_dataa_w,
		datab => add_1_datab_w,
		result => wire_altfp_div_csa8_result
	  );
	altfp_div_srt_ext1 :  Float_32_Div_altfp_div_srt_ext_14f
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		denom => man_b_w,
		divider => wire_altfp_div_srt_ext1_divider,
		numer => man_a_w,
		quotient => wire_altfp_div_srt_ext1_quotient,
		remain => wire_altfp_div_srt_ext1_remain
	  );
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_dffe <= exp_man_and_or_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_dffe1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_dffe1a <= and_or_pipeline_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_dffe3a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_dffe3a <= and_or_int_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline0c <= and_or_dffe_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline10c <= and_or_pipeline9c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline11c <= and_or_pipeline10c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline12c <= and_or_pipeline11c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline13c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline13c <= and_or_pipeline12c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline14c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline14c <= and_or_pipeline13c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline15c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline15c <= and_or_pipeline14c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline16c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline16c <= and_or_pipeline15c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline17c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline17c <= and_or_pipeline16c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline18c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline18c <= and_or_pipeline17c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline19c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline19c <= and_or_pipeline18c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline1c <= and_or_pipeline0c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline20c <= and_or_pipeline19c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline21c <= and_or_pipeline20c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline22c <= and_or_pipeline21c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline23c <= and_or_pipeline22c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline24c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline24c <= and_or_pipeline23c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline25c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline25c <= and_or_pipeline24c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline26c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline26c <= and_or_pipeline25c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline27c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline27c <= and_or_pipeline26c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline2c <= and_or_pipeline1c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline3c <= and_or_pipeline2c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline4c <= and_or_pipeline3c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline5c <= and_or_pipeline4c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline6c <= and_or_pipeline5c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline7c <= and_or_pipeline6c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline8c <= and_or_pipeline7c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN and_or_pipeline9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN and_or_pipeline9c <= and_or_pipeline8c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN bias_addition_overf_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN bias_addition_overf_dffe <= bias_addition_overf_w;
			END IF;
		END IF;
	END PROCESS;
	wire_bias_addition_overf_dffe_w_lg_q781w(0) <= bias_addition_overf_dffe AND wire_w_lg_nan_w780w(0);
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN divider_pipe1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN divider_pipe1a <= wire_altfp_div_srt_ext1_divider;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN division_by_zero_port_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN division_by_zero_port_dffe <= division_by_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_a_and_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_a_and_dffe <= exp_a_and_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_a_b_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_a_b_dffe <= exp_or_result_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_a_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_a_dffe <= wire_w_dataa_int_range365w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_a_or_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_a_or_dffe <= exp_a_or_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_a_or_dffe_w_lg_q629w(0) <= NOT exp_a_or_dffe;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_b_and_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_b_and_dffe <= exp_b_and_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_b_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_b_dffe <= wire_w_datab_int_range367w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_b_or_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_b_or_dffe <= exp_b_or_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_exp_b_or_dffe_w_lg_q632w(0) <= NOT exp_b_or_dffe;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe1a <= exp_pipeline_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_dffe2a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_dffe2a <= exp_dffe1a_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline0c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline0c <= exp_sub_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline10c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline10c <= exp_pipeline9c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline11c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline11c <= exp_pipeline10c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline12c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline12c <= exp_pipeline11c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline13c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline13c <= exp_pipeline12c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline14c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline14c <= exp_pipeline13c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline15c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline15c <= exp_pipeline14c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline16c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline16c <= exp_pipeline15c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline17c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline17c <= exp_pipeline16c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline18c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline18c <= exp_pipeline17c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline19c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline19c <= exp_pipeline18c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline1c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline1c <= exp_pipeline0c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline20c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline20c <= exp_pipeline19c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline21c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline21c <= exp_pipeline20c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline22c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline22c <= exp_pipeline21c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline23c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline23c <= exp_pipeline22c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline24c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline24c <= exp_pipeline23c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline25c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline25c <= exp_pipeline24c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline26c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline26c <= exp_pipeline25c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline2c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline2c <= exp_pipeline1c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline3c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline3c <= exp_pipeline2c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline4c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline4c <= exp_pipeline3c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline5c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline5c <= exp_pipeline4c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline6c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline6c <= exp_pipeline5c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline7c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline7c <= exp_pipeline6c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline8c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline8c <= exp_pipeline7c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_pipeline9c <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_pipeline9c <= exp_pipeline8c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN exp_res_pipe3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN exp_res_pipe3 <= exp_res_int_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN implied_bit <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN implied_bit <= wire_altfp_div_srt_ext1_quotient(26);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN implied_bit2a <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN implied_bit2a <= implied_bit;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_a_and_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_a_and_dffe <= man_a_and_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_a_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_a_dffe <= wire_w_dataa_int_range366w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_a_or_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_a_or_dffe <= man_a_or_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_man_a_or_dffe_w_lg_q635w(0) <= NOT man_a_or_dffe;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_b_and_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_b_and_dffe <= man_b_and_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_b_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_b_dffe <= wire_w_datab_int_range368w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_b_or_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_b_or_dffe <= man_b_or_msb2_w;
			END IF;
		END IF;
	END PROCESS;
	wire_man_b_or_dffe_w_lg_q638w(0) <= NOT man_b_or_dffe;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN man_res_pipe3 <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN man_res_pipe3 <= man_res_int_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN quotient_pipe1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN quotient_pipe1a <= wire_altfp_div_srt_ext1_quotient;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN remainder_pipe1a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN remainder_pipe1a <= wire_altfp_div_srt_ext1_remain;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN result_output_dffe <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN result_output_dffe <= mux_3_res_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rnd_overflow_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN rnd_overflow_dffe <= rnd_overflow;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN rnded_man_pipe2a <= (OTHERS => '0');
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN rnded_man_pipe2a <= rnded_man_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_a_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_a_dffe <= dataa_int(31);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_b_dffe <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_b_dffe <= datab_int(31);
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline0c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline0c <= sign_div;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline10c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline10c <= sign_div_pipeline9c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline11c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline11c <= sign_div_pipeline10c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline12c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline12c <= sign_div_pipeline11c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline13c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline13c <= sign_div_pipeline12c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline14c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline14c <= sign_div_pipeline13c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline15c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline15c <= sign_div_pipeline14c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline16c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline16c <= sign_div_pipeline15c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline17c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline17c <= sign_div_pipeline16c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline18c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline18c <= sign_div_pipeline17c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline19c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline19c <= sign_div_pipeline18c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline1c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline1c <= sign_div_pipeline0c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline20c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline20c <= sign_div_pipeline19c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline21c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline21c <= sign_div_pipeline20c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline22c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline22c <= sign_div_pipeline21c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline23c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline23c <= sign_div_pipeline22c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline24c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline24c <= sign_div_pipeline23c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline25c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline25c <= sign_div_pipeline24c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline26c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline26c <= sign_div_pipeline25c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline27c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline27c <= sign_div_pipeline26c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline2c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline2c <= sign_div_pipeline1c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline3c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline3c <= sign_div_pipeline2c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline4c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline4c <= sign_div_pipeline3c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline5c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline5c <= sign_div_pipeline4c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline6c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline6c <= sign_div_pipeline5c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline7c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline7c <= sign_div_pipeline6c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline8c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline8c <= sign_div_pipeline7c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_div_pipeline9c <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_div_pipeline9c <= sign_div_pipeline8c;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe1a <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe1a <= sign_div_pipeline_w;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe2a <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe2a <= sign_pipe1a;
			END IF;
		END IF;
	END PROCESS;
	PROCESS (clock, aclr)
	BEGIN
		IF (aclr = '1') THEN sign_pipe3a <= '0';
		ELSIF (clock = '1' AND clock'event) THEN 
			IF (clk_en = '1') THEN sign_pipe3a <= sign_pipe2a;
			END IF;
		END IF;
	END PROCESS;
	add_sub10 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "ADD",
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		dataa => exp_dffe2a_w,
		datab => bias_add_w,
		overflow => wire_add_sub10_overflow,
		result => wire_add_sub10_result
	  );
	add_sub9 :  lpm_add_sub
	  GENERIC MAP (
		LPM_DIRECTION => "SUB",
		LPM_PIPELINE => 1,
		LPM_REPRESENTATION => "SIGNED",
		LPM_WIDTH => 9
	  )
	  PORT MAP ( 
		aclr => aclr,
		clken => clk_en,
		clock => clock,
		dataa => exp_sub_a_w,
		datab => exp_sub_b_w,
		result => wire_add_sub9_result
	  );
	cmpr2 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 14
	  )
	  PORT MAP ( 
		aeb => wire_cmpr2_aeb,
		agb => wire_cmpr2_agb,
		dataa => quo_msb_m1_compare_dataa(52 DOWNTO 39),
		datab => quo_msb_m1_compare_datab(52 DOWNTO 39)
	  );
	cmpr3 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aeb => wire_cmpr3_aeb,
		agb => wire_cmpr3_agb,
		dataa => quo_msb_m1_compare_dataa(38 DOWNTO 26),
		datab => quo_msb_m1_compare_datab(38 DOWNTO 26)
	  );
	cmpr4 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		aeb => wire_cmpr4_aeb,
		agb => wire_cmpr4_agb,
		dataa => quo_msb_m1_compare_dataa(25 DOWNTO 13),
		datab => quo_msb_m1_compare_datab(25 DOWNTO 13)
	  );
	cmpr5 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 13
	  )
	  PORT MAP ( 
		ageb => wire_cmpr5_ageb,
		dataa => quo_msb_m1_compare_dataa(12 DOWNTO 0),
		datab => quo_msb_m1_compare_datab(12 DOWNTO 0)
	  );
	cmpr6 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 27
	  )
	  PORT MAP ( 
		aeb => wire_cmpr6_aeb,
		agb => wire_cmpr6_agb,
		dataa => quo_msb_m2_compare_dataa(53 DOWNTO 27),
		datab => quo_msb_m2_compare_datab(53 DOWNTO 27)
	  );
	cmpr7 :  lpm_compare
	  GENERIC MAP (
		LPM_REPRESENTATION => "UNSIGNED",
		LPM_WIDTH => 27
	  )
	  PORT MAP ( 
		ageb => wire_cmpr7_ageb,
		dataa => quo_msb_m2_compare_dataa(26 DOWNTO 0),
		datab => quo_msb_m2_compare_datab(26 DOWNTO 0)
	  );

 END RTL; --Float_32_Div_altfp_div_01j
--VALID FILE


LIBRARY ieee;
USE ieee.std_logic_1164.all;

ENTITY Float_32_Div IS
	PORT
	(
		clock		: IN STD_LOGIC ;
		dataa		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		datab		: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
		division_by_zero		: OUT STD_LOGIC ;
		result		: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
END Float_32_Div;


ARCHITECTURE RTL OF float_32_div IS

	SIGNAL sub_wire0	: STD_LOGIC ;
	SIGNAL sub_wire1	: STD_LOGIC_VECTOR (31 DOWNTO 0);



	COMPONENT Float_32_Div_altfp_div_01j
	PORT (
			clock	: IN STD_LOGIC ;
			dataa	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			datab	: IN STD_LOGIC_VECTOR (31 DOWNTO 0);
			division_by_zero	: OUT STD_LOGIC ;
			result	: OUT STD_LOGIC_VECTOR (31 DOWNTO 0)
	);
	END COMPONENT;

BEGIN
	division_by_zero    <= sub_wire0;
	result    <= sub_wire1(31 DOWNTO 0);

	Float_32_Div_altfp_div_01j_component : Float_32_Div_altfp_div_01j
	PORT MAP (
		clock => clock,
		dataa => dataa,
		datab => datab,
		division_by_zero => sub_wire0,
		result => sub_wire1
	);



END RTL;

-- ============================================================
-- CNX file retrieval info
-- ============================================================
-- Retrieval info: PRIVATE: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: PRIVATE: SYNTH_WRAPPER_GEN_POSTFIX STRING "0"
-- Retrieval info: LIBRARY: altera_mf altera_mf.altera_mf_components.all
-- Retrieval info: CONSTANT: DENORMAL_SUPPORT STRING "NO"
-- Retrieval info: CONSTANT: INTENDED_DEVICE_FAMILY STRING "Cyclone IV E"
-- Retrieval info: CONSTANT: OPTIMIZE STRING "AREA"
-- Retrieval info: CONSTANT: PIPELINE NUMERIC "33"
-- Retrieval info: CONSTANT: REDUCED_FUNCTIONALITY STRING "NO"
-- Retrieval info: CONSTANT: WIDTH_EXP NUMERIC "8"
-- Retrieval info: CONSTANT: WIDTH_MAN NUMERIC "23"
-- Retrieval info: USED_PORT: clock 0 0 0 0 INPUT NODEFVAL "clock"
-- Retrieval info: USED_PORT: dataa 0 0 32 0 INPUT NODEFVAL "dataa[31..0]"
-- Retrieval info: USED_PORT: datab 0 0 32 0 INPUT NODEFVAL "datab[31..0]"
-- Retrieval info: USED_PORT: division_by_zero 0 0 0 0 OUTPUT NODEFVAL "division_by_zero"
-- Retrieval info: USED_PORT: result 0 0 32 0 OUTPUT NODEFVAL "result[31..0]"
-- Retrieval info: CONNECT: @clock 0 0 0 0 clock 0 0 0 0
-- Retrieval info: CONNECT: @dataa 0 0 32 0 dataa 0 0 32 0
-- Retrieval info: CONNECT: @datab 0 0 32 0 datab 0 0 32 0
-- Retrieval info: CONNECT: division_by_zero 0 0 0 0 @division_by_zero 0 0 0 0
-- Retrieval info: CONNECT: result 0 0 32 0 @result 0 0 32 0
-- Retrieval info: GEN_FILE: TYPE_NORMAL Float_32_Div.vhd TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Float_32_Div.inc FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Float_32_Div.cmp TRUE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Float_32_Div.bsf FALSE
-- Retrieval info: GEN_FILE: TYPE_NORMAL Float_32_Div_inst.vhd TRUE
-- Retrieval info: LIB_FILE: lpm
